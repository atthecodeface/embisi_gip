/*a Copyright Gavin J Stark, 2004
 */

/*a Includes
 */
include "postbus.h"
include "gip.h"
include "io_block.h"
include "io_slots_eth_ss_par.h"
include "io_cmd.h"
include "memories.h"

/*a Types
 */

/*a External modules required
 */
/*m apb_devices
 */
extern module apb_devices( clock int_clock,
                           input bit int_reset,

                           input bit apb_pselect,
                           input bit apb_penable,
                           input bit apb_prnw,
                           input bit[6] apb_paddr,
                           input bit[32] apb_pwdata,
                           output bit[32] apb_prdata,
                           output bit apb_pwait,

                           output bit global_apb_pselect,
                           output bit global_apb_penable,
                           output bit global_apb_prnw,
                           output bit[5] global_apb_paddr,
                           output bit[32] global_apb_pwdata,
                           input bit[32] global_apb_prdata,
                           input bit global_apb_pwait,

                           output bit txd,
                           input bit rxd,

                           output bit[4]ext_bus_ce,
                           output bit ext_bus_oe,
                           output bit ext_bus_we,
                           output bit[24]ext_bus_address,
                           output bit ext_bus_write_data_enable,
                           output bit[32]ext_bus_write_data,
                           input bit[32]ext_bus_read_data,

                           input bit[4]gpio_input,
                           output bit[16]gpio_output,
                           output bit[16]gpio_output_enable,
                           output bit gpio_input_event,

                           output bit[3] timer_equalled
    )
{
    timing to rising clock int_clock int_reset;

    timing to rising clock int_clock apb_pselect, apb_penable, apb_prnw, apb_paddr, apb_pwdata;
    timing from rising clock int_clock apb_prdata, apb_pwait;

    timing from rising clock int_clock global_apb_pselect, global_apb_penable, global_apb_prnw, global_apb_paddr, global_apb_pwdata;
    timing to rising clock int_clock global_apb_prdata, global_apb_pwait;

    timing to rising clock int_clock rxd;
    timing from rising clock int_clock txd;

    timing from rising clock int_clock ext_bus_ce, ext_bus_oe, ext_bus_we, ext_bus_address, ext_bus_write_data_enable, ext_bus_write_data;
    timing to rising clock int_clock ext_bus_read_data;

    timing to rising clock int_clock gpio_input;
    timing from rising clock int_clock gpio_output, gpio_output_enable, gpio_input_event;

    timing from rising clock int_clock timer_equalled;

}

/*m gip_core_plus
 */
extern module gip_core_plus( clock int_clock,
                             input bit int_reset,

                             output bit gip_mem_priority,
                             output bit gip_mem_read,
                             output bit gip_mem_write,
                             output bit[4] gip_mem_write_byte_enables,
                             output bit[32] gip_mem_address,
                             output bit[32] gip_mem_write_data,
                             input bit[32] gip_mem_read_data,
                             input bit gip_mem_wait,

                             output bit[6] apb_paddr,
                             output bit apb_penable,
                             output bit apb_pselect,
                             output bit[32] apb_pwdata,
                             output bit apb_prnw,
                             input bit[32] apb_prdata,
                             input bit apb_pwait,

                             input bit[8] local_events_in,

                             output t_postbus_type postbus_tx_type,
                             output t_postbus_data postbus_tx_data,
                             input t_postbus_ack postbus_tx_ack,

                             input t_postbus_type postbus_rx_type,
                             input t_postbus_data postbus_rx_data,
                             output t_postbus_ack postbus_rx_ack
    )
{
    timing to rising clock int_clock int_reset;

    timing from rising clock int_clock gip_mem_priority, gip_mem_read, gip_mem_write, gip_mem_write_byte_enables, gip_mem_address, gip_mem_write_data;
    timing to rising clock int_clock gip_mem_read_data, gip_mem_wait;

    timing from rising clock int_clock apb_pselect, apb_penable, apb_prnw, apb_paddr, apb_pwdata;
    timing to rising clock int_clock apb_prdata, apb_pwait;

    timing to rising clock int_clock local_events_in;

    timing from rising clock int_clock postbus_tx_type, postbus_tx_data;
    timing to rising clock int_clock postbus_tx_ack;

    timing from rising clock int_clock postbus_rx_ack;
    timing to rising clock int_clock postbus_rx_type, postbus_rx_data;
}

/*m gip_simple_boot_rom
 */
extern module gip_simple_boot_rom( clock rom_clock,
                                   input bit rom_reset,
                                   input bit rom_read,
                                   input bit[12] rom_address,
                                   output bit[32] rom_read_data )
{
    timing to rising clock rom_clock rom_reset, rom_read, rom_address;
    timing from rising clock rom_clock rom_read_data;
}

/*m postbus_test_rom_contents
 */
extern module postbus_test_rom_contents( clock int_clock, input bit int_reset, input bit read, input bit[8] address, output bit[32] data )
{
    timing to rising clock int_clock int_reset, read, address;
    timing from rising clock int_clock data;
    timing comb input int_reset;
}

/*m ddr_dram_as_sram
 */
extern module ddr_dram_as_sram( clock drm_clock,
                                //clock slow_clock,

                                input bit drm_ctl_reset,
                                output bit init_done,

                                input bit sram_priority,
                                input bit sram_read,
                                input bit sram_write,
                                input bit[4] sram_write_byte_enables,
                                input bit[24] sram_address,
                                input bit[32] sram_write_data,
                                output bit[32] sram_read_data,
                                output bit sram_low_priority_wait,

                                input bit cke_last_of_logic,
                                output bit next_cke,
                                output bit[2] next_s_n,
                                output bit next_ras_n,
                                output bit next_cas_n,
                                output bit next_we_n,
                                output bit[13] next_a,
                                output bit[2] next_ba,
                                output bit[32] next_dq,
                                output bit[4] next_dqm,
                                output bit next_dqoe,
                                output bit[4] next_dqs_high,
                                output bit[4] next_dqs_low,
                                input bit[32] input_dq_high,
                                input bit[32] input_dq_low )
{
    timing to rising clock drm_clock cke_last_of_logic;
    timing to rising clock drm_clock drm_ctl_reset;
    timing from rising clock drm_clock init_done;

    timing from rising clock drm_clock next_cke, next_s_n, next_ras_n, next_cas_n, next_we_n, next_a, next_ba, next_dq, next_dqm, next_dqoe, next_dqs_high, next_dqs_low;
    timing to rising clock drm_clock input_dq_high, input_dq_low;

//    timing to rising clock slow_clock sram_priority, sram_read, sram_write, sram_write_byte_enables, sram_address, sram_write_data;
//    timing from rising clock slow_clock sram_read_data, sram_low_priority_wait;
}

/*m analyzer
 */
extern module analyzer( clock analyzer_clock,
                        clock output_clock,
                        clock apb_clock,

                        input bit analyzer_reset,

                        input bit[3] apb_paddr,
                        input bit apb_penable,
                        input bit apb_pselect,
                        input bit[32] apb_pwdata,
                        input bit apb_prnw,
                        output bit[32] apb_prdata,
                        output bit apb_pwait,

                        output bit trace_ready,
                        output bit trace_done,

                        output bit[32]analyzer_mux_control,
                        input bit[32]internal_signal_in,

                        input bit ext_trigger_reset,
                        input bit ext_trigger_enable,

                        input bit async_trace_read_enable,
                        output bit async_trace_valid_out,
                        output bit[32] async_trace_out )
{
    timing to rising clock analyzer_clock internal_signal_in;
    timing to rising clock analyzer_clock analyzer_reset;

    timing to rising clock output_clock ext_trigger_enable, ext_trigger_reset;
    timing to rising clock output_clock async_trace_read_enable;
    timing from rising clock output_clock async_trace_valid_out, async_trace_out;

    timing to rising clock apb_clock apb_pselect, apb_penable, apb_prnw, apb_paddr, apb_pwdata;
    timing from rising clock apb_clock apb_prdata, apb_pwait;

    timing from rising clock apb_clock trace_ready, trace_done;

}

/*a Modules
 */
module gip_system( clock drm_clock,
                   clock int_clock,
                   input bit system_reset,
                   output bit reset_out,

                   input bit[8] switches,
                   output bit[8] leds,

                   output bit txd,
                   input bit rxd,

                   output bit[4]ext_bus_ce,
                   output bit ext_bus_oe,
                   output bit ext_bus_we,
                   output bit[24]ext_bus_address,
                   output bit ext_bus_write_data_enable,
                   output bit[32]ext_bus_write_data,
                   input bit[32]ext_bus_read_data,

                   input bit cke_last_of_logic,
                   output bit next_cke,
                   output bit[2] next_s_n,
                   output bit next_ras_n,
                   output bit next_cas_n,
                   output bit next_we_n,
                   output bit[13] next_a,
                   output bit[2] next_ba,
                   output bit[32] next_dq,
                   output bit[4] next_dqm,
                   output bit next_dqoe,
                   output bit[4] next_dqs_high,
                   output bit[4] next_dqs_low,
                   input bit[32] input_dq_high,
                   input bit[32] input_dq_low,

                   clock eth_mii_tx_clock,
                   output bit eth_mii_tx_en,
                   output bit[4] eth_mii_tx_d,
                   output bit eth_mii_tx_er, // we hold this low

                   clock eth_mii_rx_clock,
                   input bit eth_mii_rx_dv,
                   input bit[4] eth_mii_rx_d,
                   input bit eth_mii_rx_er,

                   input bit eth_mii_col,
                   input bit eth_mii_crs,

                   output bit[2] sscl,
                   output bit[2] sscl_oe,
                   output bit ssdo,
                   output bit ssdo_oe,
                   input bit[2] ssdi,
                   output bit[8] sscs,

                   clock par_clock,
                   input bit[3] par_control_inputs,
                   input bit[16] par_data_inputs,

                   output bit[4] par_control_outputs,
                   output bit[4] par_control_oes,
                   output bit[16] par_data_outputs,
                   output bit[3] par_data_output_width,
                   output bit par_data_oe,

                   clock analyzer_clock,
                   output bit analyzer_async_trace_valid,
                   output bit[32] analyzer_async_trace_out
                   )
{
    default clock int_clock;
    default reset system_reset;

    comb bit int_reset;

    net bit txd;

    net bit[4]ext_bus_ce;
    net bit ext_bus_oe;
    net bit ext_bus_we;
    net bit[24]ext_bus_address;
    net bit ext_bus_write_data_enable;
    net bit[32]ext_bus_write_data;

    net bit next_cke;
    net bit[2] next_s_n;
    net bit next_ras_n;
    net bit next_cas_n;
    net bit next_we_n;
    net bit[13] next_a;
    net bit[2] next_ba;
    net bit[32] next_dq;
    net bit[4] next_dqm;
    net bit next_dqoe;
    net bit[4] next_dqs_high;
    net bit[4] next_dqs_low;

    net bit gip_mem_priority;
    net bit gip_mem_read;
    net bit gip_mem_write;
    net bit[4] gip_mem_write_byte_enables;
    net bit[32] gip_mem_address;
    net bit[32] gip_mem_write_data;
    comb bit[32] gip_mem_read_data;
    comb bit gip_mem_wait;

    net bit[6] apb_paddr;
    net bit apb_penable;
    net bit apb_pselect;
    net bit[32] apb_pwdata;
    net bit apb_prnw;
    net bit[32] apb_prdata;
    net bit apb_pwait;

    net t_postbus_type postbus_tx_type;
    net t_postbus_data postbus_tx_data;
    net t_postbus_ack postbus_tx_ack;

    net t_postbus_type postbus_rx_type;
    net t_postbus_data postbus_rx_data;
    net t_postbus_ack postbus_rx_ack;

    net bit    io_slot_cfg_write "asserted if cfg_data should be written to cfg_slot";
    net bit[8] io_slot_cfg_data  "data for setting a slot configuration";
    net bit[2] io_slot_cfg_slot  "number of slot cfg data is destined for";

    net bit[4]    io_slot_egr_cmd_ready  "bus of command emptys from all slots - they are filled asynchronously to requests";
    net bit       io_slot_egr_data_req    "OR of data requests, masked by pending acknowledgements";
    net t_io_tx_data_fifo_cmd   io_slot_egr_data_cmd    "data command from lowest number slot with an unmasked request";
    net bit[2]    io_slot_egr_data_slot   "slot the data command is coming from";
    net bit      io_slot_egr_data_ack "asserted to acknowledge the current data request";
    net bit[32]  io_slot_egr_data "contains data for writes to the slots, registered here, valid 3 cycles after acknowledged request (acked req in cycle 0, sram req in cycle 1, sram data stored end cycle 2, this valid in cycle 3";
    net bit[2]   io_slot_egr_slot "indicates which slot the egress data is for, registered here; ";
    net bit      io_slot_egr_cmd_write  "asserted if the data on the bus in this cycle is for the command side interface - if so, it will drive the not empty signal to the slot client";
    net bit      io_slot_egr_data_write "asserted if the data on the bus in this cycle is for the data side interface";

    net bit[32]  io_slot_ingr_data       "muxed in slot head from clients, ANDed with a select from io_slot_ing_number";
    net bit      io_slot_ingr_status_req "OR of status requests, masked by pending acknowledgements";
    net bit      io_slot_ingr_data_req    "OR of rx data requests, masked by pending acknowledgements, clear if status_req is asserted";
    net bit[2]   io_slot_ingr_slot       "indicates which slot the status or rx data request is from";
    net bit     io_slot_ingr_ack        "acknowledge, valid in same clock as status_req and data_req";
    net bit[4]  io_slot_ingr_data_full  "for use by I/O";

    comb bit rom_next_access;
    comb bit sram_next_access;
    comb bit dram_next_access;
    clocked bit rom_current_access = 0;
    clocked bit sram_current_access = 0;
    clocked bit dram_current_access = 0;
    net bit[32] rom_read_data;
    net bit[32] sram_read_data;
    net bit[32] dram_read_data;
    net bit dram_wait;

    net bit ddr_ready;

    comb bit io_reset;
    net bit eth_mii_tx_en;
    net bit[4] eth_mii_tx_d;
//    comb bit eth_mii_tx_er;

    net bit[16] gpio_output;
    net bit[16] gpio_output_enable;
    net bit gpio_input_event;
    net bit[3] timer_equalled;

    net bit[2] sscl;
    net bit[2] sscl_oe;
    net bit ssdo;
    net bit ssdo_oe;
    net bit[8] sscs;

    net bit[4]                par_control_outputs;
    net bit[4]                par_control_oes;
    net bit[16]               par_data_outputs;
    net bit[3]                par_data_output_width;
    net bit                   par_data_oe;

    comb bit[8] local_events_in;

    net bit[32] analyzer_mux_control;
    net bit[32] iob_analyzer_signals;
    net bit[32] ios_analyzer_signals;
    clocked bit[32] analyzer_signals = 0;
    net bit analyzer_trace_ready;
    net bit analyzer_trace_done;
    net bit analyzer_async_trace_valid;
    net bit[32] analyzer_async_trace_out;

    net bit global_apb_pselect;
    net bit global_apb_penable;
    net bit global_apb_prnw;
    net bit[5] global_apb_paddr;
    net bit[32] global_apb_pwdata;
    net bit[32] global_apb_prdata;
    net bit global_apb_pwait;

    /*b Reset detect from ethernet
      Note that the MII_RX clock stops when our reset goes off, so our reset should come from 
     */
    clocked clock eth_mii_rx_clock reset system_reset bit[8] eth_reset_count=0;
    clocked clock int_clock reset system_reset bit[3] eth_reset_shf=0;
    clocked clock int_clock reset system_reset bit eth_reset=0;
    reset_from_eth "Generate reset from incoming ethernet packet":
        {
            if (eth_mii_rx_dv && (eth_mii_rx_d==5))
            {
                eth_reset_count <= eth_reset_count+1;
            }
            else
            {
                eth_reset_count <= 0;
            }

            eth_reset_shf[0] <= (eth_reset_count[4;4]==15);
            eth_reset_shf[2;1] <= eth_reset_shf[2;0];

            eth_reset <= (eth_reset_shf[2;1]==2b01); // rising edge of eth_reset_shf synchronizer
            reset_out = system_reset || eth_reset;
        }

    /*b GIP core
     */
    gip_core "GIP core instance":
        {
            local_events_in = 0;
            local_events_in[3;0] = timer_equalled;
            local_events_in[3] = gpio_input_event;
            leds = gpio_output[8;0];
            gip_core_plus gip( int_clock <- int_clock,
                               int_reset <= int_reset,

                               gip_mem_priority => gip_mem_priority,
                               gip_mem_read => gip_mem_read,
                               gip_mem_write => gip_mem_write,
                               gip_mem_write_byte_enables => gip_mem_write_byte_enables,
                               gip_mem_address => gip_mem_address,
                               gip_mem_write_data => gip_mem_write_data,
                               gip_mem_read_data <= gip_mem_read_data,
                               gip_mem_wait <= gip_mem_wait,

                               apb_paddr => apb_paddr,
                               apb_penable => apb_penable,
                               apb_pselect => apb_pselect,
                               apb_pwdata => apb_pwdata,
                               apb_prnw => apb_prnw,
                               apb_prdata <= apb_prdata,
                               apb_pwait <= apb_pwait,

                               local_events_in <= local_events_in,

                               postbus_tx_type => postbus_tx_type,
                               postbus_tx_data => postbus_tx_data,
                               postbus_tx_ack <= postbus_tx_ack,

                               postbus_rx_type <= postbus_rx_type,
                               postbus_rx_data <= postbus_rx_data,
                               postbus_rx_ack => postbus_rx_ack );
        }

    /*b Memory subsystem
     */
    memory_subsystem "Memory subsystem":
        {
            int_reset = reset_out || !ddr_ready;

            rom_next_access = !gip_mem_address[16] && !gip_mem_address[31];
            sram_next_access = gip_mem_address[16] && !gip_mem_address[31];
            dram_next_access = !rom_next_access && !sram_next_access;
            rom_current_access <= rom_next_access;
            sram_current_access <= sram_next_access;
            dram_current_access <= dram_next_access;

            gip_simple_boot_rom boot_rom( rom_clock <- int_clock,
                                          rom_reset <= int_reset,
                                          rom_read <= rom_next_access && gip_mem_read,
                                          rom_address <= gip_mem_address[12;2],
                                          rom_read_data => rom_read_data );

            memory_s_sp_4096_x_4b8 shared_sram( sram_clock <- int_clock,
                                                sram_address <= gip_mem_address[12;2],
                                                sram_read <= sram_next_access && gip_mem_read,
                                                sram_write <= sram_next_access && gip_mem_write,
                                                sram_byte_enables <= gip_mem_write_byte_enables,
                                                sram_write_data <= gip_mem_write_data,
                                                sram_read_data => sram_read_data );

            ddr_dram_as_sram main_ram( drm_clock <- drm_clock,
                                       //slow_clock <- int_clock,

                                       drm_ctl_reset <= reset_out,
                                       init_done => ddr_ready,
                                       
                                       sram_priority <= gip_mem_priority,
                                       sram_read <= dram_next_access && gip_mem_read,
                                       sram_write <= dram_next_access && gip_mem_write,
                                       sram_write_byte_enables <= gip_mem_write_byte_enables,
                                       sram_address <= gip_mem_address[24;2],
                                       sram_write_data <= gip_mem_write_data,
                                       sram_read_data => dram_read_data,
                                       sram_low_priority_wait => dram_wait,

                                       cke_last_of_logic <= cke_last_of_logic,
                                       next_cke => next_cke,
                                       next_s_n => next_s_n,
                                       next_ras_n => next_ras_n,
                                       next_cas_n => next_cas_n,
                                       next_we_n => next_we_n,
                                       next_a => next_a,
                                       next_ba => next_ba,
                                       next_dq => next_dq,
                                       next_dqm => next_dqm,
                                       next_dqoe => next_dqoe,
                                       next_dqs_high => next_dqs_high,
                                       next_dqs_low => next_dqs_low,
                                       input_dq_high <= input_dq_high,
                                       input_dq_low <= input_dq_low );

            gip_mem_read_data = dram_read_data;
            if (rom_current_access)
            {
                gip_mem_read_data = rom_read_data;
            }
            if (sram_current_access)
            {
                gip_mem_read_data = sram_read_data;
            }
            gip_mem_wait = dram_next_access ? dram_wait : 0;

        }

    /*b APB devices
     */
    apb_devices_instanced "APB devices":
        {
            apb_devices apb( int_clock <- int_clock,
                             int_reset <= int_reset,

                             apb_pselect <= apb_pselect,
                             apb_penable <= apb_penable,
                             apb_paddr <= apb_paddr,
                             apb_prnw <= apb_prnw,
                             apb_pwdata <= apb_pwdata,
                             apb_prdata => apb_prdata,
                             apb_pwait => apb_pwait,

                             global_apb_pselect => global_apb_pselect,
                             global_apb_penable => global_apb_penable,
                             global_apb_paddr => global_apb_paddr,
                             global_apb_prnw => global_apb_prnw,
                             global_apb_pwdata => global_apb_pwdata,
                             global_apb_prdata <= global_apb_prdata,
                             global_apb_pwait <= global_apb_pwait,

                             txd => txd,
                             rxd <= rxd,

                             ext_bus_ce => ext_bus_ce,
                             ext_bus_oe => ext_bus_oe,
                             ext_bus_we => ext_bus_we,
                             ext_bus_address => ext_bus_address,
                             ext_bus_write_data_enable => ext_bus_write_data_enable,
                             ext_bus_write_data => ext_bus_write_data,
                             ext_bus_read_data <= ext_bus_read_data,
                             gpio_input <= switches[4;0],
                             gpio_output => gpio_output,
                             gpio_output_enable => gpio_output_enable,
                             gpio_input_event => gpio_input_event,

                             timer_equalled => timer_equalled
                );
        }

    /*b Postbus instances
     */
    postbus_instances "Postbus instances":
        {

            io_reset = int_reset;
            eth_mii_tx_er = 0;
            io_block iob_a( int_clock <- int_clock,
                          int_reset <= int_reset,

                          postbus_tgt_type <= postbus_tx_type,
                          postbus_tgt_data <= postbus_tx_data,
                          postbus_tgt_ack => postbus_tx_ack,

                          postbus_src_type => postbus_rx_type,
                          postbus_src_data => postbus_rx_data,
                          postbus_src_ack <= postbus_rx_ack,

                          io_slot_cfg_write => io_slot_cfg_write,
                          io_slot_cfg_data => io_slot_cfg_data,
                          io_slot_cfg_slot => io_slot_cfg_slot,

                          io_slot_egr_cmd_ready <= io_slot_egr_cmd_ready,
                          io_slot_egr_data_req <= io_slot_egr_data_req,
                            io_slot_egr_data_cmd <= io_slot_egr_data_cmd,
                          io_slot_egr_data_slot <= io_slot_egr_data_slot,
                          io_slot_egr_data_ack => io_slot_egr_data_ack,
                          io_slot_egr_data => io_slot_egr_data,
                          io_slot_egr_slot => io_slot_egr_slot,
                          io_slot_egr_cmd_write => io_slot_egr_cmd_write,
                          io_slot_egr_data_write => io_slot_egr_data_write,

                          io_slot_ingr_data <= io_slot_ingr_data,
                          io_slot_ingr_status_req <= io_slot_ingr_status_req,
                          io_slot_ingr_data_req <= io_slot_ingr_data_req,
                          io_slot_ingr_slot <= io_slot_ingr_slot,
                          io_slot_ingr_ack => io_slot_ingr_ack,
                          io_slot_ingr_data_full => io_slot_ingr_data_full,

                          analyzer_mux_control <= analyzer_mux_control[3;0],
                          analyzer_signals => iob_analyzer_signals );

            io_slots_eth_ss_par ios_a ( int_clock <- int_clock,
                                        int_reset <= int_reset,

                                        io_slot_cfg_write <= io_slot_cfg_write,
                                        io_slot_cfg_data <= io_slot_cfg_data,
                                        io_slot_cfg_slot <= io_slot_cfg_slot,

                                        io_slot_egr_cmd_ready => io_slot_egr_cmd_ready,
                                        io_slot_egr_data_req => io_slot_egr_data_req,
                                        io_slot_egr_data_cmd => io_slot_egr_data_cmd,
                                        io_slot_egr_data_slot => io_slot_egr_data_slot,
                                        io_slot_egr_data_ack <= io_slot_egr_data_ack,
                                        io_slot_egr_data <= io_slot_egr_data,
                                        io_slot_egr_slot <= io_slot_egr_slot,
                                        io_slot_egr_cmd_write <= io_slot_egr_cmd_write,
                                        io_slot_egr_data_write <= io_slot_egr_data_write,

                                        io_slot_ingr_data => io_slot_ingr_data,
                                        io_slot_ingr_status_req => io_slot_ingr_status_req,
                                        io_slot_ingr_data_req => io_slot_ingr_data_req,
                                        io_slot_ingr_slot => io_slot_ingr_slot,
                                        io_slot_ingr_ack <= io_slot_ingr_ack,
                                        io_slot_ingr_data_full <= io_slot_ingr_data_full,

                                        erx_clock <- eth_mii_rx_clock,
                                        erx_reset <= io_reset,

                                        erx_mii_dv <= eth_mii_rx_dv,
                                        erx_mii_err <= eth_mii_rx_er,
                                        erx_mii_data <= eth_mii_rx_d,

                                        etx_clock <- eth_mii_tx_clock,
                                        etx_reset <= io_reset,
                                        etx_mii_enable => eth_mii_tx_en,
                                        etx_mii_data => eth_mii_tx_d,
                                        etx_mii_crs <= eth_mii_crs,
                                        etx_mii_col <= eth_mii_col,

                                        sscl => sscl,
                                        sscl_oe => sscl_oe,
                                        ssdo => ssdo,
                                        ssdo_oe => ssdo_oe,
                                        ssdi <= ssdi,
                                        sscs => sscs,

                                        par_clock <- par_clock,
                                        par_control_inputs <= par_control_inputs,
                                        par_data_inputs <= par_data_inputs,

                                        par_control_outputs => par_control_outputs,
                                        par_control_oes => par_control_oes,
                                        par_data_outputs => par_data_outputs,
                                        par_data_output_width => par_data_output_width,
                                        par_data_oe => par_data_oe,

                                        analyzer_mux_control <= analyzer_mux_control[2;0],
                                        analyzer_signals => ios_analyzer_signals );
        }

    /*b Logic analyzer
     */
    logic_analyzer "Logic analyzer instantiation and signal muxing":
        {

            analyzer_signals <= iob_analyzer_signals;
            part_switch (analyzer_mux_control)
                {
                case 0:
                {
                    analyzer_signals <= gip_mem_address;
                    analyzer_signals[31] <= gip_mem_read;
                    analyzer_signals[30] <= gip_mem_write;
                    analyzer_signals[4;26] <= gip_mem_write_byte_enables;
                }
                case 1:
                {
                    if (gip_mem_read || gip_mem_write)
                    {
                        analyzer_signals <= gip_mem_address; // transaction type in bits [2;0] is 00->data read, 01->ins read, 10->data word write, 11->data subword write
                    }
                    else
                    {
                        analyzer_signals <= 0;
                    }
                    analyzer_signals[2;0] <= 0;
                    if (gip_mem_priority) // data read has bits 1:0 as 1
                    {
                        analyzer_signals[2;0] <= 1;
                    }
                    if (gip_mem_write) // data write (no inst write :-) has bits 1:0 as 2 or 3
                    {
                        analyzer_signals[2;0] <= 2;
                        if (gip_mem_write_byte_enables!=4hf)
                        {
                            analyzer_signals[0] <= 1;
                        }
                    }
                }
                case 4:
                {
                    analyzer_signals <= gip_mem_write_data;
                }
                case 5:
                {
                    analyzer_signals <= gip_mem_read_data;
                }
                }
            analyzer logic_analyzer( analyzer_clock <- int_clock,
                                     output_clock <- analyzer_clock,
                                     apb_clock <- int_clock,

                                     analyzer_reset <= switches[6],

                                     apb_paddr <= global_apb_paddr[3;0],
                                     apb_penable <= global_apb_penable,
                                     apb_pselect <= global_apb_pselect,
                                     apb_prnw <= global_apb_prnw,
                                     apb_pwdata <= global_apb_pwdata,
                                     apb_pwait => global_apb_pwait,
                                     apb_prdata => global_apb_prdata,

                                     trace_ready => analyzer_trace_ready,
                                     trace_done => analyzer_trace_done,

                                     analyzer_mux_control => analyzer_mux_control,
                                     internal_signal_in <= analyzer_signals,

                                     ext_trigger_reset <= 0,
                                     ext_trigger_enable <= 0,

                                     async_trace_read_enable <= switches[5],
                                     async_trace_valid_out => analyzer_async_trace_valid,
                                     async_trace_out => analyzer_async_trace_out );

        }
}

