/*a Copyright Gavin J Stark, 2004
 */

/*a To do
 */

/*a Includes
 */
include "gip.h"
include "gip_internal.h"
include "postbus.h"

/*a Constants
 */

/*a Types
 */
/*t t_gip_postbus_rx_fsm
 */
typedef fsm {
    gip_postbus_rx_fsm_idle; // Waiting for first data - go to hold or buffer_last
    gip_postbus_rx_fsm_hold; // Buffer full - write data, then go to data state
    gip_postbus_rx_fsm_data; // Buffer empty, write data directly to RF (if not GIP) and buffer in case
    gip_postbus_rx_fsm_buffer_last; // Buffer full with last word - write data
    gip_postbus_rx_fsm_signal; // All done, now just set the correct semaphore if reqd
} t_gip_postbus_rx_fsm;

/*t t_gip_postbus_tx_fsm
 */
typedef fsm
{
    gip_postbus_tx_fsm_idle; // Waiting for command pending - go to present_single or first
    gip_postbus_tx_fsm_present_single; // Single word transaction ongoing
    gip_postbus_tx_fsm_present_first; // First word of multiword transaction ongoing
    gip_postbus_tx_fsm_hold; // In the middle of a transaction, waiting for data from RF (GIP stole RF cycles)
    gip_postbus_tx_fsm_present_middle; // In the middle of a transaction presenting data
    gip_postbus_tx_fsm_present_last; // Presenting the last word of a transaction
    gip_postbus_tx_fsm_signal; // Setting the semaphore, single cycle (unless rx is setting semaphore too)
} t_gip_postbus_tx_fsm;

/*t t_gip_postbus_fifo
 */
typedef struct
{
    bit[5] base;
    bit[5] end;
    bit[5] read;
    bit[5] write;
} t_gip_postbus_fifo;

typedef struct
{
    t_gip_word a;
} t_gip_word_a;

/*a Module
 */
constant integer gip_postbus_nfifo=2;
constant integer gip_postbus_log_nfifo=1;
module gip_postbus( clock gip_clock,
                    input bit gip_reset,

                    input bit read,
                    input bit flush,
                    input bit[5] read_address,
                    output bit[32] read_data,

                    input bit write,
                    input bit[5] write_address,
                    input bit[32] write_data,

                    output t_postbus_type postbus_tx_type,
                    output t_postbus_data postbus_tx_data,
                    input t_postbus_ack postbus_tx_ack,

                    input t_postbus_type postbus_rx_type,
                    input t_postbus_data postbus_rx_data,
                    output t_postbus_ack postbus_rx_ack,

                    output bit[5] semaphore_to_set "Semaphore to set due to postbus receive/transmit - none if zero"

    )
{
    /*b Default clock and reset
     */
    default clock gip_clock;
    default reset gip_reset;

    /*b State in the special registers guaranteed by the design - note we also have a 32x32 register file, single read, single write port
     */
    net bit[32] rf_read_data;
    clocked t_gip_word_a[gip_postbus_nfifo] command = { {a=0} }; // 32-bit command registers, used in tx; includes length (in words) for transfer
    clocked t_gip_word_a[gip_postbus_nfifo] status = { {a=0} }; // 32-bit status registers, used in rx; basically user-defined data
    clocked t_gip_postbus_fifo[gip_postbus_nfifo] tx_fifo = {{base=0, end=0, read=0, write=0}}; // 4 write FIFOs - just read/write pointers, base, end, 5-bits each
    clocked t_gip_postbus_fifo[gip_postbus_nfifo] rx_fifo = {{base=0, end=0, read=0, write=0}}; // 4 read FIFOs - just read/write pointers, base, end, 5-bits each
    clocked bit[32] postbus_rx_buffer = 0; // One word store for transfer to the rf if it is being read by GIP

    clocked bit[gip_postbus_log_nfifo] postbus_rx_fifo = 0; // 0 for rx transfer to rx_fifo[0], 1 for transfer to rx_fifo[1], etc
    clocked t_gip_postbus_rx_fsm postbus_rx_fsm = gip_postbus_rx_fsm_idle; // FSM for receive side of postbus
    clocked bit postbus_rx_last = 0; // 1 if this is the first word and last word

    clocked bit[gip_postbus_nfifo] pending_tx_xfrs = 0; // 1 bit for each command, indicating transfers pending
    clocked bit[gip_postbus_log_nfifo] postbus_tx_fifo = 0; // 0 for tx transfer from tx_fifo[0], 1 for transfer from tx_fifo[1], etc
    clocked t_gip_postbus_tx_fsm postbus_tx_fsm = gip_postbus_tx_fsm_idle; // FSM for transmit side of postbus
    clocked t_postbus_data postbus_tx_data = 0; // Postbus Tx side data presented
    clocked bit[5] postbus_tx_left = 0; // Words left to transmit (0=>last)
    clocked bit[5] postbus_tx_semaphore = 0; // Semaphore to set on completion of transmit

    /*b Combinatorials in the postbus registers
     */
    comb bit[gip_postbus_log_nfifo] postbus_next_tx_fifo;

    comb bit gip_rf_write; // 1 if the GIP wants to write
    comb bit[5] gip_rf_write_r; // rf entry the GIP wants to write
    comb bit postbus_rf_write; // 1 if the postbus wants to write
    comb bit[5] postbus_rf_write_r; // rf entry the postbus wants to write
    comb bit postbus_buffer_write; // 1 if the postbus wants to write to its buffer

    comb bit gip_rf_read; // 1 if the GIP wants to read
    comb bit[5] gip_rf_read_r; // rf entry the GIP wants to read
    comb bit postbus_rf_read; // 1 if the postbus wants to read
    comb bit[5] postbus_rf_read_r; // rf entry the postbus wants to read

    comb bit clock_tx_fifo_read;
    comb bit clock_tx_fifo_write;
    comb bit clock_rx_fifo_read;
    comb bit clock_rx_fifo_write;
    comb bit tx_fifo_read_okay;
    comb bit rx_fifo_written_okay;

    comb bit[gip_postbus_log_nfifo] read_fifo;
    comb bit[gip_postbus_log_nfifo] write_fifo;

    /*b Decode the GIP request
     */
    gip_decode "Decode the GIP request":
        {
            read_fifo = read_address[gip_postbus_log_nfifo;gip_postbus_reg_fifo_bit];
            clock_rx_fifo_read = 0;
            gip_rf_read = 0;
            gip_rf_read_r = rx_fifo[read_fifo].read;
            read_data = 0;

            write_fifo = write_address[gip_postbus_log_nfifo;gip_postbus_reg_fifo_bit];
            clock_tx_fifo_write = 0;
            gip_rf_write = 0;
            gip_rf_write_r = tx_fifo[write_fifo].write;

            part_switch (read_address)
                {
                case gip_postbus_reg_status_0:
                case gip_postbus_reg_status_1:
                case gip_postbus_reg_status_2:
                case gip_postbus_reg_status_3:
                {
                    read_data[gip_postbus_nfifo;8] = pending_tx_xfrs;
                    read_data[1] = (rx_fifo[read_fifo].read != rx_fifo[read_fifo].write);
                    read_data[0] = pending_tx_xfrs[read_fifo];
                }
                case gip_postbus_reg_command_0:
                case gip_postbus_reg_command_1:
                case gip_postbus_reg_command_2:
                case gip_postbus_reg_command_3:
                {
//                    read_data = command[read_fifo].a;
                }
                case gip_postbus_reg_rx_fifo_0:
                case gip_postbus_reg_rx_fifo_1:
                case gip_postbus_reg_rx_fifo_2:
                case gip_postbus_reg_rx_fifo_3:
                {
                    if (read)
                    {
                        gip_rf_read = 1;
                        if (!flush)
                        {
                            clock_rx_fifo_read = 1;
                        }
                    }
                    read_data = rf_read_data;
                }
                case gip_postbus_reg_tx_fifo_config_0:
                case gip_postbus_reg_tx_fifo_config_1:
                case gip_postbus_reg_tx_fifo_config_2:
                case gip_postbus_reg_tx_fifo_config_3:
                {
                    read_data[5; 0] = tx_fifo[read_fifo].base;
                    read_data[5; 8] = tx_fifo[read_fifo].end;
                    read_data[5;16] = tx_fifo[read_fifo].read;
                    read_data[5;24] = tx_fifo[read_fifo].write;
                }
                case gip_postbus_reg_rx_fifo_config_0:
                case gip_postbus_reg_rx_fifo_config_1:
                case gip_postbus_reg_rx_fifo_config_2:
                case gip_postbus_reg_rx_fifo_config_3:
                {
                    read_data[5; 0] = rx_fifo[read_fifo].base;
                    read_data[5; 8] = rx_fifo[read_fifo].end;
                    read_data[5;16] = rx_fifo[read_fifo].read;
                    read_data[5;24] = rx_fifo[read_fifo].write;
                }
                }

            part_switch (write_address)
                {
                case gip_postbus_reg_command_0:
                case gip_postbus_reg_command_1:
                case gip_postbus_reg_command_2:
                case gip_postbus_reg_command_3:
                {
                    if (write)
                    {
                        command[write_fifo].a <= write_data;
                    }
                }
                case gip_postbus_reg_tx_fifo_0:
                case gip_postbus_reg_tx_fifo_1:
                case gip_postbus_reg_tx_fifo_2:
                case gip_postbus_reg_tx_fifo_3:
                {
                    if (write)
                    {
                        gip_rf_write = 1;
                        clock_tx_fifo_write = 1;
                    }
                }
                }
        }

    /*b Instantiate the RF
     */
    rf_instance "Register file instance":
        {
            rf_1r_1w_32_32 rf( rf_clock <- gip_clock,
                               rf_reset <= gip_reset,
                               rf_rd_addr_0 <= gip_rf_read ? gip_rf_read_r : postbus_rf_read_r,
                               rf_rd_data_0 => rf_read_data,
                               rf_wr_enable <= gip_rf_write | postbus_rf_write,
                               rf_wr_addr <= gip_rf_write ? gip_rf_write_r : postbus_rf_write_r,
                               rf_wr_data <= gip_rf_write ? write_data : 0  ); //postbus_rx_data of some form; register or input data
        }

    /*b Decode the FSMs
     */
    fsm_decode "Postbus FSM decodes":
        {
            semaphore_to_set = 0; // 0 means no semaphore to set
            postbus_rf_read = 0;
            postbus_rf_read_r = tx_fifo[postbus_tx_fifo].read;

            postbus_tx_type = postbus_word_type_idle;
            full_switch (postbus_tx_fsm)
                {
                case gip_postbus_tx_fsm_idle:
                {
                    postbus_tx_type = postbus_word_type_idle;
                }
                case gip_postbus_tx_fsm_present_single:
                {
                    postbus_tx_type = postbus_word_type_start;
                }
                case gip_postbus_tx_fsm_present_first:
                {
                    postbus_tx_type = postbus_word_type_start;
                    postbus_rf_read = 1;
                }
                case gip_postbus_tx_fsm_hold:
                {
                    postbus_tx_type = postbus_word_type_hold;
                    postbus_rf_read = 1;
                }
                case gip_postbus_tx_fsm_present_middle:
                {
                    postbus_tx_type = postbus_word_type_data;
                    postbus_rf_read = 1;
                }
                case gip_postbus_tx_fsm_present_last:
                {
                    postbus_tx_type = postbus_word_type_last;
                }
                case gip_postbus_tx_fsm_signal:
                {
                    postbus_tx_type = postbus_word_type_idle;
                    semaphore_to_set = postbus_tx_semaphore;
                }
                }

            postbus_rx_ack = postbus_ack_hold;
            full_switch (postbus_rx_fsm)
                {
                case gip_postbus_rx_fsm_idle:
                case gip_postbus_rx_fsm_data:
                {
                    postbus_rx_ack = postbus_ack_taken;
                }
                case gip_postbus_rx_fsm_buffer_last:
                case gip_postbus_rx_fsm_hold:
                {
                    postbus_rx_ack = postbus_ack_hold;
                }
                case gip_postbus_rx_fsm_signal:
                {
                    postbus_rx_ack = postbus_ack_hold;
//                    semaphore_to_set = status[postbus_rx_fifo].a[5;postbus_command_rx_signal_start];
                }
                }
        }

    /*b Handle FIFO pointers
     */
    fifo_pointers "Handle FIFO pointers":
        {
            if (clock_tx_fifo_read)
            {
                tx_fifo[postbus_tx_fifo].read <= tx_fifo[postbus_tx_fifo].read+1;
                if ( (tx_fifo[postbus_tx_fifo].read+1) == tx_fifo[postbus_tx_fifo].end)
                {
                    tx_fifo[postbus_tx_fifo].read <= tx_fifo[postbus_tx_fifo].base;
                }
            }
            if (clock_rx_fifo_read)
            {
                rx_fifo[read_fifo].read <= rx_fifo[read_fifo].read+1;
                if ((rx_fifo[read_fifo].read+1)==rx_fifo[read_fifo].end)
                {
                    rx_fifo[read_fifo].read <= rx_fifo[read_fifo].base;
                }
            }
            if (clock_rx_fifo_write)
            {
                rx_fifo[postbus_rx_fifo].write <= rx_fifo[postbus_rx_fifo].write+1;
                if ((rx_fifo[postbus_rx_fifo].write+1)==rx_fifo[postbus_rx_fifo].end)
                {
                    rx_fifo[postbus_rx_fifo].write <= rx_fifo[postbus_rx_fifo].base;
                }
            }
            if (clock_tx_fifo_write)
            {
                tx_fifo[write_fifo].write <= tx_fifo[write_fifo].write+1;
                if ((tx_fifo[write_fifo].write+1) == tx_fifo[write_fifo].end)
                {
                    tx_fifo[write_fifo].write <= tx_fifo[write_fifo].base;
                }
            }
            part_switch (write_address)
                {
                case gip_postbus_reg_tx_fifo_config_0:
                case gip_postbus_reg_tx_fifo_config_1:
                case gip_postbus_reg_tx_fifo_config_2:
                case gip_postbus_reg_tx_fifo_config_3:
                {
                    if (write)
                    {
                        tx_fifo[write_fifo].base  <= write_data[5; 0];
                        tx_fifo[write_fifo].end   <= write_data[5; 8];
                        tx_fifo[write_fifo].read  <= write_data[5;16];
                        tx_fifo[write_fifo].write <= write_data[5;24];
                    }
                }
                case gip_postbus_reg_rx_fifo_config_0:
                case gip_postbus_reg_rx_fifo_config_1:
                case gip_postbus_reg_rx_fifo_config_2:
                case gip_postbus_reg_rx_fifo_config_3:
                {
                    if (write)
                    {
                        rx_fifo[write_fifo].base  <= write_data[5; 0];
                        rx_fifo[write_fifo].end   <= write_data[5; 8];
                        rx_fifo[write_fifo].read  <= write_data[5;16];
                        rx_fifo[write_fifo].write <= write_data[5;24];
                    }
                }
                }
        }

    /*b Handle the Tx FSM
     */
    tx_fsm "Postbus transmit FSM":
        {
            clock_tx_fifo_read = 0;
            tx_fifo_read_okay = !gip_rf_read;
            postbus_next_tx_fifo = 0;
            full_switch (postbus_tx_fsm)
            {
            case gip_postbus_tx_fsm_idle:
            {
                if (pending_tx_xfrs!=0)
                {
                    full_switch (pending_tx_xfrs)
                        {
                        case 1:
                        case 3:
                        case 5:
                        case 7:
                        case 9:
                        case 4hb:
                        case 4hd:
                        case 4hf:
                        {
                            postbus_next_tx_fifo = 0;
                        }
                        case 2:
                        case 6:
                        case 4ha:
                        case 4he:
                        {
                            postbus_next_tx_fifo = 1;
                        }
                        case 4:
                        case 4hc:
                        {
                            postbus_next_tx_fifo = 2;
                        }
                        case 8:
                        {
                            postbus_next_tx_fifo = 3;
                        }
                        }

                    postbus_tx_data <= command[ postbus_next_tx_fifo ].a;
                    postbus_tx_semaphore <= command[postbus_next_tx_fifo].a[5;postbus_command_tx_signal_start];
                    if (command[ postbus_next_tx_fifo ].a[postbus_command_last_bit])
                    {
                        postbus_tx_fsm <= gip_postbus_tx_fsm_present_single;
                    }
                    else
                    {
                        postbus_tx_fsm <= gip_postbus_tx_fsm_present_first;
                    }
                    postbus_tx_left <= command[ postbus_next_tx_fifo ].a[5;postbus_command_tx_length_start];
                    postbus_tx_fifo <= postbus_next_tx_fifo;
                }
            }
            case gip_postbus_tx_fsm_present_single:
            {
                if (postbus_tx_ack == postbus_ack_taken)
                {
                    postbus_tx_fsm <= gip_postbus_tx_fsm_signal;
                }
            }
            case gip_postbus_tx_fsm_present_first:
            case gip_postbus_tx_fsm_present_middle: 
            {
                if (postbus_tx_ack == postbus_ack_taken)
                {
                    if (tx_fifo_read_okay)
                    {
                        clock_tx_fifo_read = 1; // move on FIFO ptr, decrement length
                        if (postbus_tx_left == 0)
                        {
                            postbus_tx_fsm <= gip_postbus_tx_fsm_present_last;
                        }
                        else
                        {
                            postbus_tx_fsm <= gip_postbus_tx_fsm_present_middle;
                        }
                    }
                    else
                    {
                        postbus_tx_fsm <= gip_postbus_tx_fsm_hold;
                    }
                }
                else
                {
                    postbus_tx_fsm <= postbus_tx_fsm; // Making it clear this is okay for both single and middle
                }
            }
            case gip_postbus_tx_fsm_hold:
            {
                if (tx_fifo_read_okay)
                {
                    clock_tx_fifo_read = 1; // move on FIFO ptr, decrement length
                    if (postbus_tx_left == 0)
                    {
                        postbus_tx_fsm <= gip_postbus_tx_fsm_present_last;
                    }
                    else
                    {
                        postbus_tx_fsm <= gip_postbus_tx_fsm_present_middle;
                    }
                }
            }
            case gip_postbus_tx_fsm_present_last:
            {
                if (postbus_tx_ack == postbus_ack_taken)
                {
                    postbus_tx_fsm <= gip_postbus_tx_fsm_signal;
                }
            }
            case gip_postbus_tx_fsm_signal:
            {
                if (postbus_rx_fsm != gip_postbus_rx_fsm_signal)
                {
                    pending_tx_xfrs[postbus_tx_fifo] <= 0;
                    postbus_tx_fsm <= gip_postbus_tx_fsm_idle;
                }
            }
            }
            if (clock_tx_fifo_read)
            {
                postbus_tx_left <= postbus_tx_left-1;
                postbus_tx_data <= rf_read_data;
            }
            part_switch (write_address)
                {
                case gip_postbus_reg_command_0:
                case gip_postbus_reg_command_1:
                case gip_postbus_reg_command_2:
                case gip_postbus_reg_command_3:
                {
                    if (write)
                    {
                        pending_tx_xfrs[write_fifo] <= 1;
                    }
                }
                }
        }

    /*b Handle the Rx FSM
     */
    rx_fsm "Postbus receive FSM":
        {
            postbus_rf_write = 0;
            postbus_rf_write_r = rx_fifo[0].write;
            rx_fifo_written_okay = !gip_rf_write;
            postbus_buffer_write = 0;
            full_switch (postbus_rx_fsm)
            {
            case gip_postbus_rx_fsm_idle:
            {
                if (postbus_rx_type != postbus_word_type_idle)
                {
                    postbus_rx_fsm <= gip_postbus_rx_fsm_hold;
                    postbus_rx_last <= postbus_rx_data[postbus_command_last_bit];
                    postbus_buffer_write = 1;
                    postbus_rx_fifo <= postbus_rx_data[31];
                }
            }
            case gip_postbus_rx_fsm_hold:
            {
                postbus_rf_write = 1;
                if (rx_fifo_written_okay)
                {
                    if (postbus_rx_last)
                    {
                        postbus_rx_fsm <= gip_postbus_rx_fsm_signal;
                    }
                    else
                    {
                        postbus_rx_fsm <= gip_postbus_rx_fsm_data;
                    }
                }
            }
            case gip_postbus_rx_fsm_data:
            {
                postbus_buffer_write = 1;
                postbus_rf_write = 1;
                postbus_rx_last <= 0;
                part_switch (postbus_rx_type)
                {
                case postbus_word_type_data:
                case postbus_word_type_start: // we treat start as data - its defensive
                {
                    if (!rx_fifo_written_okay)
                    {
                        postbus_rx_fsm <= gip_postbus_rx_fsm_hold;
                    }
                }
                case postbus_word_type_last:
                {
                    if (rx_fifo_written_okay)
                    {
                        postbus_rx_fsm <= gip_postbus_rx_fsm_signal;
                    }
                    else
                    {
                        postbus_rx_fsm <= gip_postbus_rx_fsm_buffer_last;
                    }
                }
                }
            }
            case gip_postbus_rx_fsm_buffer_last:
            {
                postbus_rf_write = 1;
                if (rx_fifo_written_okay)
                {
                    postbus_rx_fsm <= gip_postbus_rx_fsm_signal;
                }
            }
            case gip_postbus_rx_fsm_signal:
            {
                postbus_rx_last <= 0;
                postbus_rx_fsm <= gip_postbus_rx_fsm_idle; // We assume the signalling always works
            }
            }
            clock_rx_fifo_write = 0;
            if (postbus_buffer_write)
            {
                postbus_rx_buffer <= postbus_rx_data;
                clock_rx_fifo_write = rx_fifo_written_okay;
            }
        }

    /*b Done
     */
}
