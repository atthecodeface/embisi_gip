/*a To do
  Reduce gate count
  make ldm and stm use CP for non-zero cycles
 */

/*a Includes
 */
include "gip.h"
include "gip_internal.h"
include "arm.h"

/*a Types
 */

/*a Module
 */
module gip_decode_arm( input bit[32] opcode,
                       input bit[5] cycle_of_opcode,

                       output t_gip_instruction_rf inst,
                       output bit arm_use_native_decode,

                       output bit[5] next_cycle_of_opcode,
                       output t_gip_pc_op pc_op,
                       output bit[32] arm_branch_offset,

                       input bit extended,
                       input bit[28] extended_immediate,
                       input t_gip_ins_r extended_rd,
                       input t_gip_ins_r extended_rn,
                       input t_gip_ins_r extended_rm,
                       input t_gip_ext_cmd extended_cmd,

                       input bit[16] stored_reg_set,
                       output bit[16] next_stored_reg_set
                       )
{
    comb bit[4] cc;
    comb bit conditional;
    comb bit[4] alu_op;
    comb bit alu_sign;
    comb bit alu_imm;

    comb bit rd_is_pc;

    comb bit[4] alu_imm_rotate;
    comb bit[8] alu_imm_val;
    comb bit[32] alu_immediate;
    comb bit[4] alu_rd;
    comb bit[4] alu_rn;
    comb bit[4] alu_rm;
    comb bit[4] alu_rs;

    comb bit[5] alu_shf_imm_amt;
    comb bit[2] alu_shf_how;
    comb bit alu_shf_by_reg;
    comb bit alu_lsl_by_imm_0;

    comb bit ld_st_imm;
    comb bit ld_st_pre;
    comb bit ld_st_up;
    comb bit ld_st_byte;
    comb bit ld_st_wb;
    comb bit[12] ld_st_offset;

    comb bit[16] ldm_stm_reg_set;
    comb bit[5] ldm_stm_num_regs;
    comb bit[16] sel_reg_set;
    comb bit[4] ldm_stm_bottom_bit_set;

    comb t_gip_ins_cc ins_cc;
    comb t_gip_ins_cc inv_cc;

    comb t_gip_ins_r arm_mapped_rn;
    comb t_gip_ins_r arm_mapped_rd;
    comb t_gip_ins_r arm_mapped_rm;
    comb t_gip_ins_r arm_mapped_rs;
    comb t_gip_ins_r arm_mapped_bottom_bit_set;

    comb t_arm_ins_class ins_class;

    comb t_gip_ins_class alu_gip_ins_class;
    comb t_gip_ins_subclass alu_gip_ins_subclass;
    comb t_gip_ins_subclass alu_gip_shf;
    comb bit alu_gip_set_acc;
    comb bit alu_gip_set_flags;
    comb bit alu_gip_pass_p;
    comb bit alu_gip_set_rd;

    comb t_gip_ins_subclass ld_st_gip_ins_subclass;
    comb t_gip_ins_subclass ld_st_gip_ins_subclass_not_pre_not_post;
    comb t_gip_ins_subclass ld_st_gip_ins_subclass_post;
    comb t_gip_ins_subclass ldm_stm_gip_ins_subclass;

    comb bit branch_link;

    /*b Break out instruction and map to internal instructions
     */
    breakout_instruction "Breakout instruction":
        {
            /*b Break out the opcode
             */
            cc = opcode[4;28];
            conditional = (cc!=14);

            /*b  Break out bits for a branch
             */
            branch_link = opcode[24];
            arm_branch_offset = 0;
            arm_branch_offset[24;2] = opcode[24;0];
            if (opcode[23])
            {
                arm_branch_offset[6;26] = -1;
            }

            /*b  Break out bits for an ALU operation branch
             */
            alu_imm = opcode[25];
            alu_op = opcode[4;21];
            alu_sign = opcode[20];
            alu_imm_rotate = opcode[4;8];
            alu_imm_val = opcode[8;0];
            alu_immediate = 0;
            full_switch (alu_imm_rotate)
                {
                case 0:  { alu_immediate[8;0] = alu_imm_val; }
                case 1:  { alu_immediate[2;30] = alu_imm_val[2;0]; alu_immediate[6;0] = alu_imm_val[6;2]; }
                case 2:  { alu_immediate[4;28] = alu_imm_val[4;0]; alu_immediate[4;0] = alu_imm_val[4;4]; }
                case 3:  { alu_immediate[6;26] = alu_imm_val[6;0]; alu_immediate[2;0] = alu_imm_val[2;6]; }
                case 4:  { alu_immediate[8;24] = alu_imm_val; }
                case 5:  { alu_immediate[8;22] = alu_imm_val; }
                case 6:  { alu_immediate[8;20] = alu_imm_val; }
                case 7:  { alu_immediate[8;18] = alu_imm_val; }
                case 8:  { alu_immediate[8;16] = alu_imm_val; }
                case 9:  { alu_immediate[8;14] = alu_imm_val; }
                case 10: { alu_immediate[8;12] = alu_imm_val; }
                case 11: { alu_immediate[8;10] = alu_imm_val; }
                case 12: { alu_immediate[8;8] = alu_imm_val; }
                case 13: { alu_immediate[8;6] = alu_imm_val; }
                case 14: { alu_immediate[8;4] = alu_imm_val; }
                case 15: { alu_immediate[8;2] = alu_imm_val; }
                }

            /*b Registers
             */
            alu_rn = opcode[4;16]; // and loads/stores, ldm/stm - destination for multiplies!
            alu_rd = opcode[4;12]; // and loads/stores - rn for multiplies
            alu_rs = opcode[4;8];
            alu_rm = opcode[4;0];

            /*b Shift operation
             */
            alu_shf_imm_amt = opcode[5;7];
            alu_shf_how = opcode[2;5];
            alu_shf_by_reg = opcode[4];
            alu_lsl_by_imm_0 = 0;
            if ((alu_shf_how == arm_shf_lsl) &&
                (!alu_shf_by_reg) &&
                (alu_shf_imm_amt==0) )
            {
                alu_lsl_by_imm_0 = 1;
            }

            /*b Load/store data
             */
            ld_st_imm = !opcode[25];
            ld_st_pre = opcode[24]; // also ldm/stm
            ld_st_up = opcode[23]; // also ldm/stm
            ld_st_byte = opcode[22]; // psr in ldm/stm
            ld_st_wb = opcode[21]; // also in ldm/stm
            ld_st_offset = opcode[12;0];

            /*b LDM/STM
             */
            ldm_stm_reg_set = opcode[16;0];
            ldm_stm_num_regs = 0;
            full_switch (ldm_stm_reg_set[4;0])
                {
                case 0: {ldm_stm_num_regs = ldm_stm_num_regs+0;}
                case 1:
                case 2:
                case 4:
                case 8: {ldm_stm_num_regs = ldm_stm_num_regs+1;}
                case 3:
                case 5:
                case 6:
                case 9:
                case 10:
                case 12: {ldm_stm_num_regs = ldm_stm_num_regs+2;}
                case 7:
                case 11:
                case 13:
                case 14: {ldm_stm_num_regs = ldm_stm_num_regs+3;}
                case 15: {ldm_stm_num_regs = ldm_stm_num_regs+4;}
                }
            full_switch (ldm_stm_reg_set[4;4])
                {
                case 0: {ldm_stm_num_regs = ldm_stm_num_regs+0;}
                case 1:
                case 2:
                case 4:
                case 8: {ldm_stm_num_regs = ldm_stm_num_regs+1;}
                case 3:
                case 5:
                case 6:
                case 9:
                case 10:
                case 12: {ldm_stm_num_regs = ldm_stm_num_regs+2;}
                case 7:
                case 11:
                case 13:
                case 14: {ldm_stm_num_regs = ldm_stm_num_regs+3;}
                case 15: {ldm_stm_num_regs = ldm_stm_num_regs+4;}
                }
            full_switch (ldm_stm_reg_set[4;8])
                {
                case 0: {ldm_stm_num_regs = ldm_stm_num_regs+0;}
                case 1:
                case 2:
                case 4:
                case 8: {ldm_stm_num_regs = ldm_stm_num_regs+1;}
                case 3:
                case 5:
                case 6:
                case 9:
                case 10:
                case 12: {ldm_stm_num_regs = ldm_stm_num_regs+2;}
                case 7:
                case 11:
                case 13:
                case 14: {ldm_stm_num_regs = ldm_stm_num_regs+3;}
                case 15: {ldm_stm_num_regs = ldm_stm_num_regs+4;}
                }
            full_switch (ldm_stm_reg_set[4;12])
                {
                case 0: {ldm_stm_num_regs = ldm_stm_num_regs+0;}
                case 1:
                case 2:
                case 4:
                case 8: {ldm_stm_num_regs = ldm_stm_num_regs+1;}
                case 3:
                case 5:
                case 6:
                case 9:
                case 10:
                case 12: {ldm_stm_num_regs = ldm_stm_num_regs+2;}
                case 7:
                case 11:
                case 13:
                case 14: {ldm_stm_num_regs = ldm_stm_num_regs+3;}
                case 15: {ldm_stm_num_regs = ldm_stm_num_regs+4;}
                }
            if (cycle_of_opcode[4]==0)
            {
                sel_reg_set = ldm_stm_reg_set;
            }
            else
            {
                sel_reg_set = stored_reg_set;
            }
            ldm_stm_bottom_bit_set = 0;
            if (sel_reg_set[15]) {ldm_stm_bottom_bit_set=15;}
            if (sel_reg_set[14]) {ldm_stm_bottom_bit_set=14;}
            if (sel_reg_set[13]) {ldm_stm_bottom_bit_set=13;}
            if (sel_reg_set[12]) {ldm_stm_bottom_bit_set=12;}
            if (sel_reg_set[11]) {ldm_stm_bottom_bit_set=11;}
            if (sel_reg_set[10]) {ldm_stm_bottom_bit_set=10;}
            if (sel_reg_set[ 9]) {ldm_stm_bottom_bit_set= 9;}
            if (sel_reg_set[ 8]) {ldm_stm_bottom_bit_set= 8;}
            if (sel_reg_set[ 7]) {ldm_stm_bottom_bit_set= 7;}
            if (sel_reg_set[ 6]) {ldm_stm_bottom_bit_set= 6;}
            if (sel_reg_set[ 5]) {ldm_stm_bottom_bit_set= 5;}
            if (sel_reg_set[ 4]) {ldm_stm_bottom_bit_set= 4;}
            if (sel_reg_set[ 3]) {ldm_stm_bottom_bit_set= 3;}
            if (sel_reg_set[ 2]) {ldm_stm_bottom_bit_set= 2;}
            if (sel_reg_set[ 1]) {ldm_stm_bottom_bit_set= 1;}
            if (sel_reg_set[ 0]) {ldm_stm_bottom_bit_set= 0;}
        }

    /*b Map registers and immediate
     */
    map_registers "Map registers and immediate value using the extended amounts in the current registers (from previous instruction decodes)":
        {
            /*b Map condition code
             */
            full_switch( cc )
                {
                case 0: { ins_cc = gip_ins_cc_eq; inv_cc = gip_ins_cc_ne; }
                case 1: { ins_cc = gip_ins_cc_ne; inv_cc = gip_ins_cc_eq; }
                case 2: { ins_cc = gip_ins_cc_cs; inv_cc = gip_ins_cc_cc; }
                case 3: { ins_cc = gip_ins_cc_cc; inv_cc = gip_ins_cc_cs; }
                case 4: { ins_cc = gip_ins_cc_mi; inv_cc = gip_ins_cc_pl; }
                case 5: { ins_cc = gip_ins_cc_pl; inv_cc = gip_ins_cc_mi; }
                case 6: { ins_cc = gip_ins_cc_vs; inv_cc = gip_ins_cc_vc; }
                case 7: { ins_cc = gip_ins_cc_vc; inv_cc = gip_ins_cc_vs; }
                case 8: { ins_cc = gip_ins_cc_hi; inv_cc = gip_ins_cc_ls; }
                case 9: { ins_cc = gip_ins_cc_ls; inv_cc = gip_ins_cc_hi; }
                case 10: { ins_cc = gip_ins_cc_ge; inv_cc = gip_ins_cc_lt; }
                case 11: { ins_cc = gip_ins_cc_lt; inv_cc = gip_ins_cc_ge; }
                case 12: { ins_cc = gip_ins_cc_gt; inv_cc = gip_ins_cc_le; }
                case 13: { ins_cc = gip_ins_cc_le; inv_cc = gip_ins_cc_gt; }
                case 14: { ins_cc = gip_ins_cc_always; inv_cc = gip_ins_cc_always; }
                case 15: { ins_cc = gip_ins_cc_always; inv_cc = gip_ins_cc_always; }
                }

            /*b Map operation and setting flags
             */
//            arm_mapped_rn = map_source_register( rn );
//            arm_mapped_rm = map_source_register( shf_rm );
//            arm_mapped_rs = map_source_register( shf_rs );
//            arm_mapped_rd = map_destination_register( rd );

            /*b Map rd to instruction rd; pc if that is 15; but if extended, to full given extension
             */
            rd_is_pc = 0;
            arm_mapped_rd.type = gip_ins_r_type_register;
            arm_mapped_rd.r = 0;
            arm_mapped_rd.r[4;0] = alu_rd;
            if (alu_rd==15) { arm_mapped_rd = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc}; rd_is_pc = 1;}
            if (extended_rd.type!=gip_ins_r_type_no_override) { arm_mapped_rd = extended_rd; rd_is_pc = 0; }

            /*b Map rn to instruction rn; acc if that is 15; but if extended, to full given extension
             */
            arm_mapped_rn.type = gip_ins_r_type_register;
            arm_mapped_rn.r = 0;
            arm_mapped_rn.r[4;0] = alu_rn;
            if (alu_rn==15) { arm_mapped_rn = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc}; } // differs from native - should native match?
            if (extended_rn.type!=gip_ins_r_type_no_override) {
                arm_mapped_rn.type = extended_rn.type;
                arm_mapped_rn.r[4] = extended_rn.r[4];
                arm_mapped_rn.r[4;0] = alu_rn;
            }

            /*b Map rm to instruction rm; pc if that is 15; but if extended, to full given extension
             */
            arm_mapped_rm.type = gip_ins_r_type_register;
            arm_mapped_rm.r = 0;
            arm_mapped_rm.r[4;0] = alu_rm;
            if (alu_rm==15) { arm_mapped_rm = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc}; } // Differs from native
            if (extended_rm.type!=gip_ins_r_type_no_override)
            {
                arm_mapped_rm.type = extended_rm.type;
                arm_mapped_rm.r[4]=extended_rm.r[4];
                arm_mapped_rm.r[4;0]=alu_rm;
            }

            /*b Map rs to instruction rs; always the specified register (no extensions, PC not allowed)
             */
            arm_mapped_rs.type = gip_ins_r_type_register;
            arm_mapped_rs.r = 0;
            arm_mapped_rs.r[4;0] = alu_rs;

            /*b Map bottom bit set reg to instruction reg; no extenstions, PC allowed
             */
            arm_mapped_bottom_bit_set.type = gip_ins_r_type_register;
            arm_mapped_bottom_bit_set.r = 0;
            arm_mapped_bottom_bit_set.r[4;0] = ldm_stm_bottom_bit_set;
            if (ldm_stm_bottom_bit_set==15) { arm_mapped_bottom_bit_set = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc}; }
        }

    /*b Decode instruction class
     */
    decode_instruction_class "Decode instruction class":
        {
            ins_class = arm_ins_class_none;
            full_switch (opcode[3;25])
                {
                case 0:
                {
                    if ( (opcode[3;22]==0) &&
                         (opcode[4;4]==9) )
                    {
                        ins_class = arm_ins_class_mul;
                    }
                    else
                    {
                        ins_class = arm_ins_class_alu;
                    }
                }
                case 1:
                {
                    ins_class = arm_ins_class_alu;
                }
                case 2:
                case 3:
                {
                    if (opcode[20])
                    {
                        ins_class = arm_ins_class_load; // note also that [25] must not be 1 at the same time as a [4] being one - this is a shift by register, which is not permitted, and may be decoded as something else?
                    }
                    else
                    {
                        ins_class = arm_ins_class_store;
                    }
                }
                case 4:
                {
                    if (opcode[20])
                    {
                        ins_class = arm_ins_class_ldm;
                    }
                    else
                    {
                        ins_class = arm_ins_class_stm;
                    }
                }
                case 5:
                {
                    ins_class = arm_ins_class_branch;
                }
                case 6:
                {
                    ins_class = arm_ins_class_native;
                }
                default:
                {
                    ins_class = arm_ins_class_none;
                }
                }
        }

    /*b ARM ALU decode
     */
    arm_alu_decode "ALU instructions map to one or more internal instructions
                    Those that do not set the PC and are immediate or have a shift of LSL #0 map to one internal ALU instruction
                    Those that do not set the PC and have a shift other than LSL #0 map to one internal SHIFT instruction and one internal ALU instruction
                    Those that set the PC and have a shift of LSL #0 map to one internal ALU instruction with 'flush' set
                    Those that set the PC and have a shift other than LSL #0 map to one internal SHIFT instruction and one internal ALU instruction with 'flush' set" :
        {
            /*b Map shift type
             */
            alu_gip_shf = gip_ins_subclass_shift_lsl;
            full_switch (alu_shf_how)
                {
                case arm_shf_lsl:
                {
                    alu_gip_shf = gip_ins_subclass_shift_lsl;
                }
                case arm_shf_lsr:
                {
                    alu_gip_shf = gip_ins_subclass_shift_lsr;
                }
                case arm_shf_asr:
                {
                    alu_gip_shf = gip_ins_subclass_shift_asr;
                }
                case arm_shf_ror:
                {
                    alu_gip_shf = gip_ins_subclass_shift_ror;
                    if (!alu_shf_by_reg && (alu_shf_imm_amt==0))
                    {
                        alu_gip_shf = gip_ins_subclass_shift_ror33;
                    }
                }
                }

            /*b Map to internal GIP ALU instruction type
             */
            alu_gip_ins_class = gip_ins_class_arith;
            alu_gip_ins_subclass = gip_ins_subclass_arith_add;
            alu_gip_set_acc = 0;
            alu_gip_set_flags = 0;
            alu_gip_pass_p = 0;
            alu_gip_set_rd = 1;

            full_switch (alu_op)
                {
                case  0: // and
                {
                    alu_gip_ins_class = gip_ins_class_logic;
                    alu_gip_ins_subclass = gip_ins_subclass_logic_and;
                    alu_gip_set_flags = alu_sign;
                    alu_gip_pass_p = alu_sign;
                    alu_gip_set_acc = !conditional;
                }
                case  1: // eor
                {
                    alu_gip_ins_class = gip_ins_class_logic;
                    alu_gip_ins_subclass = gip_ins_subclass_logic_xor;
                    alu_gip_set_flags = alu_sign;
                    alu_gip_pass_p = alu_sign;
                    alu_gip_set_acc = !conditional;
                }
                case  2: // sub
                {
                    alu_gip_ins_class = gip_ins_class_arith;
                    alu_gip_ins_subclass = gip_ins_subclass_arith_sub;
                    alu_gip_set_flags = alu_sign;
                    alu_gip_set_acc = !conditional;
                }
                case  3: // rsb
                {
                    alu_gip_ins_class = gip_ins_class_arith;
                    alu_gip_ins_subclass = gip_ins_subclass_arith_rsb;
                    alu_gip_set_flags = alu_sign;
                    alu_gip_set_acc = !conditional;
                }
                case  4: // add
                {
                    alu_gip_ins_class = gip_ins_class_arith;
                    alu_gip_ins_subclass = gip_ins_subclass_arith_add;
                    alu_gip_set_flags = alu_sign;
                    alu_gip_set_acc = !conditional;
                }
                case  5: // adc
                {
                    alu_gip_ins_class = gip_ins_class_arith;
                    alu_gip_ins_subclass = gip_ins_subclass_arith_adc;
                    alu_gip_set_flags = alu_sign;
                    alu_gip_set_acc = !conditional;
                }
                case  6: // sbc
                {
                    alu_gip_ins_class = gip_ins_class_arith;
                    alu_gip_ins_subclass = gip_ins_subclass_arith_sbc;
                    alu_gip_set_flags = alu_sign;
                    alu_gip_set_acc = !conditional;
                }
                case  7: // rsc
                {
                    alu_gip_ins_class = gip_ins_class_arith;
                    alu_gip_ins_subclass = gip_ins_subclass_arith_rsc;
                    alu_gip_set_flags = alu_sign;
                    alu_gip_set_acc = !conditional;
                }
                case  8: // tst
                {
                    alu_gip_ins_class = gip_ins_class_logic;
                    alu_gip_ins_subclass = gip_ins_subclass_logic_and;
                    alu_gip_set_flags = 1;
                    alu_gip_pass_p = alu_sign;
                    alu_gip_set_acc = 0;
                    alu_gip_set_rd = 0;
                }
                case  9: // teq
                {
                    alu_gip_ins_class = gip_ins_class_logic;
                    alu_gip_ins_subclass = gip_ins_subclass_logic_xor;
                    alu_gip_set_flags = 1;
                    alu_gip_pass_p = alu_sign;
                    alu_gip_set_acc = 0;
                    alu_gip_set_rd = 0;
                }
                case 10: // cmp
                {
                    alu_gip_ins_class = gip_ins_class_arith;
                    alu_gip_ins_subclass = gip_ins_subclass_arith_sub;
                    alu_gip_set_flags = 1;
                    alu_gip_set_acc = 0;
                    alu_gip_set_rd = 0;
                }
                case 11: // cmn
                {
                    alu_gip_ins_class = gip_ins_class_arith;
                    alu_gip_ins_subclass = gip_ins_subclass_arith_add;
                    alu_gip_set_flags = 1;
                    alu_gip_set_acc = 0;
                    alu_gip_set_rd = 0;
                }
                case 12: // orr
                {
                    alu_gip_ins_class = gip_ins_class_logic;
                    alu_gip_ins_subclass = gip_ins_subclass_logic_or;
                    alu_gip_set_flags = alu_sign;
                    alu_gip_pass_p = alu_sign;
                    alu_gip_set_acc = !conditional;
                }
                case 13: // mov
                {
                    alu_gip_ins_class = gip_ins_class_logic;
                    alu_gip_ins_subclass = gip_ins_subclass_logic_mov;
                    alu_gip_set_flags = alu_sign;
                    alu_gip_pass_p = alu_sign;
                    alu_gip_set_acc = !conditional;
                }
                case 14: // bic
                {
                    alu_gip_ins_class = gip_ins_class_logic;
                    alu_gip_ins_subclass = gip_ins_subclass_logic_bic;
                    alu_gip_set_flags = alu_sign;
                    alu_gip_pass_p = alu_sign;
                    alu_gip_set_acc = !conditional;
                }
                case 15: // mvn
                {
                    alu_gip_ins_class = gip_ins_class_logic;
                    alu_gip_ins_subclass = gip_ins_subclass_logic_mvn;
                    alu_gip_set_flags = alu_sign;
                    alu_gip_pass_p = alu_sign;
                    alu_gip_set_acc = !conditional;
                }
                }
        }


    /*b Load/store decode
     */
    load_store_decode "ARM Load/store decode":
        {
            ld_st_gip_ins_subclass_not_pre_not_post = 0;
            if (ld_st_byte)
            {
                ld_st_gip_ins_subclass_not_pre_not_post = ld_st_gip_ins_subclass_not_pre_not_post | gip_ins_subclass_memory_byte;
            }
            else
            {
                ld_st_gip_ins_subclass_not_pre_not_post = ld_st_gip_ins_subclass_not_pre_not_post | gip_ins_subclass_memory_word;
            }
            if (ld_st_up)
            {
                ld_st_gip_ins_subclass_not_pre_not_post = ld_st_gip_ins_subclass_not_pre_not_post | gip_ins_subclass_memory_up;
            }
            else
            {
                ld_st_gip_ins_subclass_not_pre_not_post = ld_st_gip_ins_subclass_not_pre_not_post | gip_ins_subclass_memory_down;
            }
            ld_st_gip_ins_subclass_post = ld_st_gip_ins_subclass_not_pre_not_post | gip_ins_subclass_memory_postindex;
            if (ld_st_pre)
            {
                ld_st_gip_ins_subclass = ld_st_gip_ins_subclass_not_pre_not_post | gip_ins_subclass_memory_preindex;
            }
            else
            {
                ld_st_gip_ins_subclass = ld_st_gip_ins_subclass_not_pre_not_post | gip_ins_subclass_memory_postindex;
            }
            ldm_stm_gip_ins_subclass = gip_ins_subclass_memory_word | gip_ins_subclass_memory_up;
            if (ld_st_pre^ld_st_up)
            {
                ldm_stm_gip_ins_subclass = ldm_stm_gip_ins_subclass | gip_ins_subclass_memory_postindex;
            }
            else
            {
                ldm_stm_gip_ins_subclass = ldm_stm_gip_ins_subclass | gip_ins_subclass_memory_preindex;
            }
                                                      
        }

    /*b Decode instruction
     */
    decode_instruction "Decode instruction":
        {
            /*b Define outputs as a NOP
             */
            next_cycle_of_opcode = 0;
            pc_op = gip_pc_op_sequential;

            inst.gip_ins_class = gip_ins_class_logic;
            inst.gip_ins_subclass = gip_ins_subclass_logic_mov;
            inst.gip_ins_cc = ins_cc;
            inst.a = 0;
            inst.s_or_stack = 0;
            inst.p_or_offset_is_shift = 0;
            inst.k = 0;
            inst.f = 0;
            inst.d = 0;
            inst.gip_ins_rm = arm_mapped_rm;
            inst.gip_ins_rn = arm_mapped_rn;
            inst.gip_ins_rd = {type=gip_ins_r_type_none, r=arm_mapped_rd.r};
            inst.rm_is_imm = 0;
            inst.immediate = alu_immediate;
            inst.valid = 0;
            next_stored_reg_set = sel_reg_set;
            arm_use_native_decode = 0;

            /*b Decode instruction according to class
             */
            full_switch (ins_class)
                {
                /*b None
                 */
                case arm_ins_class_none:
                {
                    inst.valid = 0;
                }
                /*b ALU
                 */
                case arm_ins_class_alu:
                {
                    /*b Test for shift of 'LSL #0' or plain immediate
                     */
                    if (alu_imm)
                    {
                        inst.gip_ins_class =  alu_gip_ins_class;
                        inst.gip_ins_subclass =  alu_gip_ins_subclass;
                        inst.a = alu_gip_set_acc;
                        inst.s_or_stack = alu_gip_set_flags;
                        inst.p_or_offset_is_shift = 0;
                        inst.gip_ins_rm = arm_mapped_rm;
                        inst.gip_ins_rn = arm_mapped_rn;
                        inst.gip_ins_rd = arm_mapped_rd;
                        if (!alu_gip_set_rd)
                        {
                            inst.gip_ins_rd.type = gip_ins_r_type_none;
                        }
                        inst.rm_is_imm = 1;
                        inst.immediate = alu_immediate;
                        inst.valid = 1;
                        next_cycle_of_opcode = 0;
                        pc_op = gip_pc_op_sequential;
                    }
                    elsif ( alu_lsl_by_imm_0 )
                    {
                        inst.gip_ins_class =  alu_gip_ins_class;
                        inst.gip_ins_subclass =  alu_gip_ins_subclass;
                        inst.a = alu_gip_set_acc;
                        inst.s_or_stack = alu_gip_set_flags;
                        inst.p_or_offset_is_shift = 0;
                        inst.gip_ins_rm = arm_mapped_rm;
                        inst.gip_ins_rn = arm_mapped_rn;
                        inst.gip_ins_rd = arm_mapped_rd;
                        if (!alu_gip_set_rd)
                        {
                            inst.gip_ins_rd.type = gip_ins_r_type_none;
                        }
                        inst.rm_is_imm = 0;
                        inst.immediate = alu_immediate;
                        inst.valid = 1;
                        next_cycle_of_opcode = 0;
                        pc_op = gip_pc_op_sequential;
                    }
                    else
                    {
                        full_switch (cycle_of_opcode)
                        {
                        case 0:
                        {
                            inst.gip_ins_class = gip_ins_class_shift;
                            inst.gip_ins_subclass = alu_gip_shf;
                            // First one could be done always, or conditional - it does not effect flags; we do conditional
                            inst.a = 0;
                            inst.s_or_stack = 0;
                            inst.p_or_offset_is_shift = 0;
                            inst.gip_ins_rn = arm_mapped_rm; // Yes, rm
                            inst.gip_ins_rd.type = gip_ins_r_type_none;
                            inst.valid = 1;
                            if (!alu_shf_by_reg) // Immediate shift, non-zero or non-LSL: ISHF{CC} Rm, #imm; IALU{CC}(SP|)[A][F] Rn, SHF -> Rd
                            {
                                inst.rm_is_imm = 1;
                                inst.immediate = 0;
                                inst.immediate[5;0] = alu_shf_imm_amt;
                                if (alu_shf_imm_amt==0)
                                {
                                    inst.immediate[5] = 1;
                                }
                            }
                            else // if (shf_by_reg) - must be! ISHF{CC} Rm, Rs; IALU{CC}(SP|)[A][F] Rn, SHF -> Rd
                            {
                                inst.rm_is_imm = 0;
                                inst.gip_ins_rm = arm_mapped_rs;
                            }

                            inst.valid = 1;
                            next_cycle_of_opcode = 1;
                            pc_op = gip_pc_op_hold;
                        }
                        default:
                        {
                            inst.gip_ins_class =  alu_gip_ins_class;
                            inst.gip_ins_subclass =  alu_gip_ins_subclass;
                            inst.gip_ins_cc = gip_ins_cc_cp;

                            inst.a = alu_gip_set_acc;
                            inst.s_or_stack = alu_gip_set_flags;
                            inst.p_or_offset_is_shift = alu_gip_pass_p;
                            inst.gip_ins_rm = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_shf };
                            inst.gip_ins_rn = arm_mapped_rn;
                            inst.gip_ins_rd = arm_mapped_rd;
                            if (!alu_gip_set_rd)
                            {
                                inst.gip_ins_rd.type = gip_ins_r_type_none;
                            }

                            inst.valid = 1;
                            next_cycle_of_opcode = 0;
                            pc_op = gip_pc_op_sequential;
                        }
                        }
                    }
                    inst.f = 0; // Now sort out the flush - always flush if writing to the PC, never otherwise
                    if ( (inst.gip_ins_rd.type==gip_ins_r_type_internal) &&
                         (inst.gip_ins_rd.r==gip_ins_r_int_pc) )
                    {
                        inst.f = 1;
                    }
                }
                /*b Load
                 */
                case arm_ins_class_load:
                {
                    /*b Handle immediate or reg without shift - 3 cases: preindexed without writeback (maps to ILDR), preindex with writeback (maps to IADD/SUB and ILDR), or postindexed (maps to ILDR, MOV)
                     */
                    if (ld_st_imm || alu_lsl_by_imm_0) // offset with immediate or unshifted register
                    {
                        /*b Preindexed, no writeback
                         */
                        if (ld_st_pre && !ld_st_wb) // preindexed immediate/reg: ILDR[CC]A[F] #0 (Rn, #+/-imm or +/-Rm) -> Rd
                        {
                            inst.gip_ins_class = gip_ins_class_load;
                            inst.gip_ins_subclass = ld_st_gip_ins_subclass;
                            inst.a = 1;
                            inst.s_or_stack = (alu_rn==13);
                            inst.p_or_offset_is_shift = 0;

                            inst.gip_ins_rm = arm_mapped_rm;
                            inst.gip_ins_rd = arm_mapped_rd;
                            inst.gip_ins_rn = arm_mapped_rn;
                            if (ld_st_imm)
                            {
                                inst.rm_is_imm = 1;
                                inst.immediate = 0;
                                inst.immediate[12;0] = ld_st_offset;
                            }
                            else
                            {
                                inst.rm_is_imm = 0;
                            }

                            inst.f = rd_is_pc;

                            inst.valid = 1;
                            next_cycle_of_opcode = 0;
                            pc_op = gip_pc_op_sequential;
                        }
                        /*b Preindexed, writeback
                         */
                        elsif (ld_st_pre) // preindexed immediate/reg with writeback: IADD[CC]A/ISUB[CC]A Rn, #imm/Rm -> Rn; ILDRCP[F] #0, (Acc) -> Rd
                        {
                            full_switch (cycle_of_opcode)
                            {
                            case 0:
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = ld_st_up ? gip_ins_subclass_arith_add : gip_ins_subclass_arith_sub;
                                inst.a = 1;
                                inst.s_or_stack = 0;
                                inst.p_or_offset_is_shift = 0;
                                inst.gip_ins_rd = arm_mapped_rn; // writeback address register
                                inst.gip_ins_rn = arm_mapped_rn;
                                if (ld_st_imm)
                                {
                                    inst.rm_is_imm = 1;
                                    inst.immediate = 0;
                                    inst.immediate[12;0] = ld_st_offset;
                                }
                                else
                                {
                                    inst.rm_is_imm = 0;
                                }
                                inst.valid = 1;
                                next_cycle_of_opcode = 1;
                                pc_op = gip_pc_op_hold;
                            }
                            default:
                            {
                                inst.gip_ins_class = gip_ins_class_load;
                                inst.gip_ins_subclass = ld_st_gip_ins_subclass;
                                inst.gip_ins_cc = gip_ins_cc_cp;
                                inst.a = 0;
                                inst.s_or_stack = (alu_rn==13);
                                inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_acc};
                                inst.gip_ins_rd = arm_mapped_rd;
                                inst.rm_is_imm = 1;
                                inst.immediate = 0;

                                inst.f = rd_is_pc;

                                inst.valid = 1;
                                next_cycle_of_opcode = 0;
                                pc_op = gip_pc_op_sequential;
                            }
                            }
                        }
                        /*b Postindexed
                         */
                        else // postindexed immediate/reg: ILDR[CC]A #0, (Rn), +/-Rm/Imm -> Rd; MOVCP[F] Acc -> Rn
                        {
                            full_switch (cycle_of_opcode)
                            {
                            case 0:
                            {
                                inst.gip_ins_class = gip_ins_class_load;
                                inst.gip_ins_subclass = ld_st_gip_ins_subclass;
                                inst.a = 1;
                                inst.s_or_stack = (alu_rn==13);
                                inst.p_or_offset_is_shift = 0;

                                inst.gip_ins_rm = arm_mapped_rm;
                                inst.gip_ins_rd = arm_mapped_rd;
                                inst.gip_ins_rn = arm_mapped_rn;
                                if (ld_st_imm)
                                {
                                    inst.rm_is_imm = 1;
                                    inst.immediate = 0;
                                    inst.immediate[12;0] = ld_st_offset;
                                }
                                else
                                {
                                    inst.rm_is_imm = 0;
                                }
                                inst.valid = 1;
                                next_cycle_of_opcode = 1;
                                pc_op = gip_pc_op_hold;
                            }
                            default:
                            {
                                inst.gip_ins_class = gip_ins_class_logic;
                                inst.gip_ins_subclass = gip_ins_subclass_logic_mov;
                                inst.gip_ins_cc = gip_ins_cc_cp;
                                inst.a = 0;
                                inst.s_or_stack = 0;
                                inst.p_or_offset_is_shift = 0;
                                inst.gip_ins_rd = arm_mapped_rn; // writeback address register
                                inst.rm_is_imm = 0;
                                inst.gip_ins_rm = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_acc};

                                inst.f = rd_is_pc;

                                inst.valid = 1;
                                next_cycle_of_opcode = 0;
                                pc_op = gip_pc_op_sequential;
                            }
                            }
                        }
                    }
                    /*b Register with shift
                     */
                    else // reg with shift
                    {
                        /*b Preindexed without writeback
                         */
                        if (ld_st_pre && !ld_st_wb) // preindexed reg with shift: ISHF[CC] Rm, #imm; ILDRCPA[F] (Rn, +/-SHF) -> Rd
                        {
                            full_switch (cycle_of_opcode)
                            {
                            case 0:
                            {
                                inst.gip_ins_class = gip_ins_class_shift;
                                inst.gip_ins_subclass = alu_gip_shf;
                                inst.a = 0;
                                inst.s_or_stack = 0;
                                inst.p_or_offset_is_shift = 0;
                                inst.gip_ins_rn = arm_mapped_rm; // Yes, rm
                                inst.gip_ins_rd.type = gip_ins_r_type_none;
                                inst.valid = 1;

                                inst.rm_is_imm = 1;
                                inst.immediate = 0;
                                inst.immediate[5;0] = alu_shf_imm_amt;
                                if (alu_shf_imm_amt==0)
                                {
                                    inst.immediate[5] = 1;
                                }
                                inst.valid = 1;
                                next_cycle_of_opcode = 1;
                                pc_op = gip_pc_op_hold;
                            }
                            default:
                            {
                                inst.gip_ins_class = gip_ins_class_load;
                                inst.gip_ins_subclass = ld_st_gip_ins_subclass;
                                inst.gip_ins_cc = gip_ins_cc_cp;
                                inst.a = 1;
                                inst.s_or_stack = (alu_rn==13);
                                inst.gip_ins_rn = arm_mapped_rn;
                                inst.gip_ins_rd = arm_mapped_rd;
                                inst.gip_ins_rm = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_shf};
                                inst.rm_is_imm = 0;

                                inst.f = rd_is_pc;

                                inst.valid = 1;
                                next_cycle_of_opcode = 0;
                                pc_op = gip_pc_op_sequential;
                            }
                            }
                        }
                        /*b Preindexed with writeback
                         */
                        elsif (ld_st_pre) // preindexed reg with shift with writeback: ISHF[CC] Rm, #imm; IADDCPA/ISUBCPA Rn, SHF -> Rn; ILDRCP[F] #0 (Acc) -> Rd
                        {
                            full_switch (cycle_of_opcode)
                            {
                            case 0:
                            {
                                inst.gip_ins_class = gip_ins_class_shift;
                                inst.gip_ins_subclass = alu_gip_shf;
                                inst.a = 0;
                                inst.s_or_stack = 0;
                                inst.p_or_offset_is_shift = 0;
                                inst.gip_ins_rn = arm_mapped_rm; // Yes, rm
                                inst.gip_ins_rd.type = gip_ins_r_type_none;
                                inst.valid = 1;

                                inst.rm_is_imm = 1;
                                inst.immediate = 0;
                                inst.immediate[5;0] = alu_shf_imm_amt;
                                if (alu_shf_imm_amt==0)
                                {
                                    inst.immediate[5] = 1;
                                }
                                inst.valid = 1;
                                next_cycle_of_opcode = 1;
                                pc_op = gip_pc_op_hold;
                            }
                            case 1:
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = ld_st_up ? gip_ins_subclass_arith_add : gip_ins_subclass_arith_sub;
                                inst.gip_ins_cc = gip_ins_cc_cp;
                                inst.a = 1;
                                inst.s_or_stack = 0;
                                inst.p_or_offset_is_shift = 0;
                                inst.gip_ins_rd = arm_mapped_rn; // writeback address register
                                inst.gip_ins_rn = arm_mapped_rn;
                                inst.gip_ins_rm = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_shf};
                                inst.rm_is_imm = 0;
                                inst.valid = 1;
                                next_cycle_of_opcode = 2;
                                pc_op = gip_pc_op_hold;
                            }
                            default:
                            {
                                inst.gip_ins_class = gip_ins_class_load;
                                inst.gip_ins_subclass = ld_st_gip_ins_subclass;
                                inst.gip_ins_cc = gip_ins_cc_cp;
                                inst.a = 0;
                                inst.s_or_stack = (alu_rn==13);
                                inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_acc};
                                inst.gip_ins_rd = arm_mapped_rd;
                                inst.rm_is_imm = 1;
                                inst.immediate = 0;

                                inst.f = rd_is_pc;

                                inst.valid = 1;
                                next_cycle_of_opcode = 0;
                                pc_op = gip_pc_op_sequential;
                            }
                            }
                        }
                        /*b Postindexed
                         */
                        else // postindexed reg with shift with writeback: ISHF[CC] Rm, #imm; ILDRCPA #0 (Rn), +/-SHF -> Rd; MOVCP[F] Acc -> Rn
                        {
                            full_switch (cycle_of_opcode)
                            {
                            case 0:
                            {
                                inst.gip_ins_class = gip_ins_class_shift;
                                inst.gip_ins_subclass = alu_gip_shf;
                                inst.a = 0;
                                inst.s_or_stack = 0;
                                inst.p_or_offset_is_shift = 0;
                                inst.gip_ins_rn = arm_mapped_rm; // Yes, rm
                                inst.gip_ins_rd.type = gip_ins_r_type_none;
                                inst.valid = 1;

                                inst.rm_is_imm = 1;
                                inst.immediate = 0;
                                inst.immediate[5;0] = alu_shf_imm_amt;
                                if (alu_shf_imm_amt==0)
                                {
                                    inst.immediate[5] = 1;
                                }
                                inst.valid = 1;
                                next_cycle_of_opcode = 1;
                                pc_op = gip_pc_op_hold;
                            }
                            case 1:
                            {
                                inst.gip_ins_class = gip_ins_class_load;
                                inst.gip_ins_subclass = ld_st_gip_ins_subclass;
                                inst.gip_ins_cc = gip_ins_cc_cp;
                                inst.a = 1;
                                inst.s_or_stack = (alu_rn==13);
                                inst.gip_ins_rn = arm_mapped_rn;
                                inst.gip_ins_rd = arm_mapped_rd;
                                inst.gip_ins_rm = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_shf};
                                inst.rm_is_imm = 0;

                                inst.valid = 1;
                                next_cycle_of_opcode = 2;
                                pc_op = gip_pc_op_hold;

                            }
                            default:
                            {
                                inst.gip_ins_class = gip_ins_class_logic;
                                inst.gip_ins_subclass = gip_ins_subclass_logic_mov;
                                inst.gip_ins_cc = gip_ins_cc_cp;
                                inst.a = 0;
                                inst.s_or_stack = 0;
                                inst.p_or_offset_is_shift = 0;
                                inst.gip_ins_rd = arm_mapped_rn; // writeback address register
                                inst.rm_is_imm = 0;
                                inst.gip_ins_rm = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_acc};

                                inst.f = rd_is_pc;

                                inst.valid = 1;
                                next_cycle_of_opcode = 0;
                                pc_op = gip_pc_op_sequential;
                            }
                            }
                        }
                    }

                }
                /*b Store - no offset, preindexed immediate, preindexed reg, preindexed reg with shift, postindexed immediate, postindexed reg, postindexed reg with shift
                 */
                case arm_ins_class_store:
                {
                    /*b Immediate offset of zero
                     */
                    if ( ld_st_imm && (ld_st_offset==0) ) // no offset (hence no writeback, none needed); ISTR[CC] #0 (Rn) <- Rd
                    {
                        inst.gip_ins_class = gip_ins_class_store;
                        inst.gip_ins_subclass = ld_st_gip_ins_subclass_post; // Guaranteed postindex, so we don't care what the offset is
                        inst.a = 0;
                        inst.s_or_stack = (alu_rn==13);
                        inst.p_or_offset_is_shift = 0; // with postindex means we don't care what we add; we don't store accumulator anyway

                        inst.gip_ins_rm = arm_mapped_rd;
                        inst.gip_ins_rd = {type=gip_ins_r_type_none};
                        inst.gip_ins_rn = arm_mapped_rn;

                        inst.valid = 1;
                        next_cycle_of_opcode = 0;
                        pc_op = gip_pc_op_sequential;
                    }
                    /*b Preindexed store
                     */
                    elsif (ld_st_pre)
                        {
                            /*b preindexed immediate or rm no shift: IADD[CC]AC/ISUB[CC]AC Rn, #imm/Rm; ISTRCPA[S] #0, (ACC, +/-SHF) <- Rd [-> Rn]
                             */
                            if ( ld_st_imm || alu_lsl_by_imm_0 )
                            {
                                full_switch (cycle_of_opcode)
                                    {
                                    case 0: // Ensure SHF gets cleared!
                                    {
                                        inst.gip_ins_class = gip_ins_class_arith;
                                        inst.gip_ins_subclass = ld_st_up ? gip_ins_subclass_arith_add : gip_ins_subclass_arith_sub;
                                        inst.a = 1;
                                        inst.s_or_stack = 0;
                                        inst.p_or_offset_is_shift = 0;
                                        inst.gip_ins_rd = {type=gip_ins_r_type_none};
                                        inst.gip_ins_rn = arm_mapped_rn;
                                        if (ld_st_imm)
                                        {
                                            inst.rm_is_imm = 1;
                                            inst.immediate = 0;
                                            inst.immediate[12;0] = ld_st_offset;
                                        }
                                        else
                                        {
                                            inst.rm_is_imm = 0;
                                        }
                                        inst.valid = 1;
                                        next_cycle_of_opcode = 1;
                                        pc_op = gip_pc_op_hold;
                                    }
                                    default:
                                    {
                                        inst.gip_ins_class = gip_ins_class_store;
                                        inst.gip_ins_subclass = ld_st_gip_ins_subclass;
                                        inst.gip_ins_cc = gip_ins_cc_cp;
                                        inst.a = 1;
                                        inst.s_or_stack = (alu_rn==13);
                                        inst.p_or_offset_is_shift = 1;

                                        inst.gip_ins_rm = arm_mapped_rd;
                                        inst.gip_ins_rd = {type=gip_ins_r_type_none};
                                        if (ld_st_wb)
                                        {
                                            inst.gip_ins_rd = arm_mapped_rn;
                                        }
                                        inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_acc};

                                        inst.valid = 1;
                                        next_cycle_of_opcode = 0;
                                        pc_op = gip_pc_op_sequential;
                                    }
                                    }
                            }
                            /*b Preindexed Rm with shift: ISHF[CC] Rm, #imm; ISTRCPA[S] #0, (Rn, +/-SHF) <- Rd [-> Rn]
                             */
                            else
                            {
                                full_switch (cycle_of_opcode)
                                    {
                                    case 0:
                                    {
                                        inst.gip_ins_class = gip_ins_class_shift;
                                        inst.gip_ins_subclass = alu_gip_shf;
                                        inst.a = 0;
                                        inst.s_or_stack = 0;
                                        inst.p_or_offset_is_shift = 0;
                                        inst.gip_ins_rn = arm_mapped_rm; // Yes, rm
                                        inst.gip_ins_rd = {type=gip_ins_r_type_none};
                                        inst.valid = 1;

                                        inst.rm_is_imm = 1;
                                        inst.immediate = 0;
                                        inst.immediate[5;0] = alu_shf_imm_amt;
                                        if (alu_shf_imm_amt==0)
                                        {
                                            inst.immediate[5] = 1;
                                        }

                                        inst.valid = 1;

                                        next_cycle_of_opcode = 1;
                                        pc_op = gip_pc_op_hold;
                                    }
                                    default:
                                    {
                                        inst.gip_ins_class = gip_ins_class_store;
                                        inst.gip_ins_subclass = ld_st_gip_ins_subclass;
                                        inst.gip_ins_cc = gip_ins_cc_cp;
                                        inst.a = 1;
                                        inst.s_or_stack = (alu_rn==13);
                                        inst.p_or_offset_is_shift = 1;

                                        inst.gip_ins_rm = arm_mapped_rd;
                                        inst.gip_ins_rd = {type=gip_ins_r_type_none};
                                        if (ld_st_wb)
                                        {
                                            inst.gip_ins_rd = arm_mapped_rn;
                                        }
                                        inst.gip_ins_rn = arm_mapped_rn;

                                        inst.valid = 1;

                                        next_cycle_of_opcode = 0;
                                        pc_op = gip_pc_op_sequential;
                                    }
                                    }
                            }
                        }
                    /*b Postindexed
                     */
                    else // if (!pre) - must be postindexed:
                    {
                        /*b Postindexed immediate or reg without shift;  ISTR[CC][S] #0 (Rn) <-Rd; IADDCPA/ISUBCPA Rn, #Imm/Rm -> Rn
                         */
                        if ( ld_st_imm || alu_lsl_by_imm_0 )
                        {
                            full_switch (cycle_of_opcode)
                                {
                                case 0:
                                {
                                    inst.gip_ins_class = gip_ins_class_store;
                                    inst.gip_ins_subclass = ld_st_gip_ins_subclass_post; // Guaranteed postindex, so we don't care what the offset is
                                    inst.a = 0;
                                    inst.s_or_stack = (alu_rn==13);
                                    inst.p_or_offset_is_shift = 0; // with postindex means we don't care what we add; we don't store accumulator anyway

                                    inst.gip_ins_rm = arm_mapped_rd;
                                    inst.gip_ins_rd = {type=gip_ins_r_type_none};
                                    inst.gip_ins_rn = arm_mapped_rn;

                                    inst.valid = 1;
                                    next_cycle_of_opcode = 1;
                                    pc_op = gip_pc_op_hold;
                                }
                                default:
                                {
                                    inst.gip_ins_class = gip_ins_class_arith;
                                    inst.gip_ins_subclass = ld_st_up ? gip_ins_subclass_arith_add : gip_ins_subclass_arith_sub;
                                    inst.gip_ins_cc = gip_ins_cc_cp;
                                    inst.a = 1;
                                    inst.s_or_stack = 0;
                                    inst.p_or_offset_is_shift = 0;
                                    inst.gip_ins_rd = arm_mapped_rn;
                                    inst.gip_ins_rn = arm_mapped_rn;
                                    if (ld_st_imm)
                                    {
                                        inst.rm_is_imm = 1;
                                        inst.immediate = 0;
                                        inst.immediate[12;0] = ld_st_offset;
                                    }
                                    else
                                    {
                                        inst.rm_is_imm = 0;
                                    }

                                    inst.valid = 1;

                                    next_cycle_of_opcode = 0;
                                    pc_op = gip_pc_op_sequential;
                                }
                                }
                        }
                        /*b Postindexed reg with shift
                         */
                        else //  ISHF[CC] Rm, #imm; ISTRCPA[S] #0 (Rn), +/-SHF) <-Rd -> Rn
                        {
                            full_switch (cycle_of_opcode)
                                {
                                case 0:
                                {
                                    inst.gip_ins_class = gip_ins_class_shift;
                                    inst.gip_ins_subclass = alu_gip_shf;
                                    inst.a = 0;
                                    inst.s_or_stack = 0;
                                    inst.p_or_offset_is_shift = 0;
                                    inst.gip_ins_rn = arm_mapped_rm; // Yes, rm
                                    inst.gip_ins_rd = {type=gip_ins_r_type_none};
                                    inst.valid = 1;

                                    inst.rm_is_imm = 1;
                                    inst.immediate = 0;
                                    inst.immediate[5;0] = alu_shf_imm_amt;
                                    if (alu_shf_imm_amt==0)
                                    {
                                        inst.immediate[5] = 1;
                                    }

                                    inst.valid = 1;

                                    next_cycle_of_opcode = 1;
                                    pc_op = gip_pc_op_hold;

                                }
                                default:
                                {
                                    inst.gip_ins_class = gip_ins_class_store;
                                    inst.gip_ins_subclass = ld_st_gip_ins_subclass;
                                    inst.gip_ins_cc = gip_ins_cc_cp;
                                    inst.a = 1;
                                    inst.s_or_stack = (alu_rn==13);
                                    inst.p_or_offset_is_shift = 1;

                                    inst.gip_ins_rm = arm_mapped_rd;
                                    inst.gip_ins_rd = {type=gip_ins_r_type_none};
                                    if (ld_st_wb)
                                    {
                                        inst.gip_ins_rd = arm_mapped_rn;
                                    }
                                    inst.gip_ins_rn = arm_mapped_rn;

                                    inst.valid = 1;

                                    next_cycle_of_opcode = 0;
                                    pc_op = gip_pc_op_sequential;
                                }
                                }
                        }
                    }
                }
                /*b Load multiple
                 */
                case arm_ins_class_ldm:
                {

                    /*b Handle first cycle, or others
                     */
                    full_switch (cycle_of_opcode)
                    {
                    case 0:
                    {
                        /*b If DB/DA, do first instruction to generate base address: ISUB[CC]A Rn, #num_regs*4 [-> Rn]
                         */
                        if (!ld_st_up)
                        {
                            inst.gip_ins_class = gip_ins_class_arith;
                            inst.gip_ins_subclass = gip_ins_subclass_arith_sub;
                            inst.a = 1;
                            inst.s_or_stack = 0;
                            inst.p_or_offset_is_shift = 0;

                            inst.gip_ins_rd = {type=gip_ins_r_type_none};
                            if (ld_st_wb)
                            {
                                inst.gip_ins_rd = arm_mapped_rn;
                            }
                            inst.gip_ins_rn = arm_mapped_rn;

                            inst.rm_is_imm = 1;
                            inst.immediate = 0;
                            inst.immediate[5;2] = ldm_stm_num_regs;

                            inst.valid = 1;

                            next_cycle_of_opcode[5;0] = ldm_stm_num_regs-1;
                            next_cycle_of_opcode[4] = 1;
                            pc_op = gip_pc_op_hold;
                        }
                        /*b Else generate a 'ILDR[CC]A[S][F] #i Rn, #+4 [->Rn] or preindexed version
                         */
                        else
                        {
                            inst.gip_ins_class = gip_ins_class_load;
                            inst.gip_ins_subclass = ldm_stm_gip_ins_subclass;
                            inst.a = 1;
                            inst.s_or_stack = (alu_rn==13);
                            inst.p_or_offset_is_shift = 0;

                            inst.gip_ins_rd = arm_mapped_bottom_bit_set;
                            inst.gip_ins_rn = arm_mapped_rn;
                            inst.k = ldm_stm_num_regs[4;0]-1;
                            inst.rm_is_imm = 1;
                            inst.immediate = 4;

                            inst.valid = 1;

                            if (ldm_stm_num_regs==1)
                            {
                                if (ld_st_wb)
                                {
                                    next_cycle_of_opcode = 1;
                                    pc_op = gip_pc_op_hold;
                                }
                                else
                                {
                                    inst.f = opcode[15];
                                    next_cycle_of_opcode = 0;
                                    pc_op = gip_pc_op_sequential;
                                }
                            }
                            else
                            {
                                next_cycle_of_opcode[5;0] = ldm_stm_num_regs-2;
                                next_cycle_of_opcode[4] = 1;
                                pc_op = gip_pc_op_hold;
                            }

                            next_stored_reg_set[ldm_stm_bottom_bit_set] = 0;

                        }
                    }
                    /*b If IB/IA with writeback then do final MOVCP[F] Acc -> Rn; F if PC was read in the list
                     */
                    case 1:
                    {
                        inst.gip_ins_class = gip_ins_class_logic;
                        inst.gip_ins_subclass = gip_ins_subclass_logic_mov;
                        inst.gip_ins_cc = gip_ins_cc_cp;
                        inst.a = 0;
                        inst.s_or_stack = 0;
                        inst.p_or_offset_is_shift = 0;
                        inst.gip_ins_rd = arm_mapped_rn; // writeback address register
                        inst.rm_is_imm = 0;
                        inst.gip_ins_rm = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_acc};

                        inst.f = opcode[15];

                        inst.valid = 1;
                        next_cycle_of_opcode = 0;
                        pc_op = gip_pc_op_sequential;
                    }
                    /*b Handle intermediate cycles - generate a 'ILDRCPA[S][F] #i (Acc), #+4 -> reg or preindexed version
                     */
                    default:
                    {
                        inst.gip_ins_class = gip_ins_class_load;
                        inst.gip_ins_subclass = ldm_stm_gip_ins_subclass;
                        inst.gip_ins_cc = gip_ins_cc_cp;
                        inst.a = 1;
                        inst.s_or_stack = (alu_rn==13);
                        inst.p_or_offset_is_shift = 0;

                        inst.gip_ins_rd = arm_mapped_bottom_bit_set;
                        inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_acc};

                        inst.rm_is_imm = 1;
                        inst.immediate = 4;

                        inst.k = cycle_of_opcode[4;0];

                        inst.valid = 1;

                        if (cycle_of_opcode[4;0]==0) // No more to do after this one
                        {
                            if (ld_st_up && ld_st_wb)
                            {
                                next_cycle_of_opcode = 1;
                                pc_op = gip_pc_op_hold;
                            }
                            else
                            {
                                if (opcode[15])
                                {
                                    inst.f = 1;
                                }
                                next_cycle_of_opcode = 0;
                                pc_op = gip_pc_op_sequential;
                            }
                        }
                        else
                        {
                            next_cycle_of_opcode[4] = 1;
                            next_cycle_of_opcode[4;0] = cycle_of_opcode[4;0]-1;
                            pc_op = gip_pc_op_hold;
                        }

                        next_stored_reg_set[ldm_stm_bottom_bit_set] = 0;

                    }
                    }

                    /*b However, if there are no registers in the original list, just ditch everything
                     */
                    if (ldm_stm_num_regs==0)
                    {
                        inst.valid = 0;
                        next_cycle_of_opcode = 0;
                        pc_op = gip_pc_op_sequential;
                    }
                }
                /*b Store multiple
                 */
                case arm_ins_class_stm:
                {
                    /*b Handle first cycle, or others
                     */
                    if (cycle_of_opcode==0)
                    {
                        /*b If DB/DA, do first instruction to generate base address: ISUB[CC]A Rn, #num_regs*4 [-> Rn]
                         */
                        if (!ld_st_up)
                        {
                            inst.gip_ins_class = gip_ins_class_arith;
                            inst.gip_ins_subclass = gip_ins_subclass_arith_sub;
                            inst.a = 1;
                            inst.s_or_stack = 0;
                            inst.p_or_offset_is_shift = 0;

                            inst.gip_ins_rd = {type=gip_ins_r_type_none};
                            if (ld_st_wb)
                            {
                                inst.gip_ins_rd = arm_mapped_rn;
                            }
                            inst.gip_ins_rn = arm_mapped_rn;

                            inst.rm_is_imm = 1;
                            inst.immediate = 0;
                            inst.immediate[5;2] = ldm_stm_num_regs;

                            inst.valid = 1;

                            next_cycle_of_opcode[5;0] = ldm_stm_num_regs-1;
                            next_cycle_of_opcode[4] = 1;
                            pc_op = gip_pc_op_hold;
                        }
                        /*b Else generate a 'ISTR[CC]A[S][F] #i Rn, #+4 [->Rn] or preindexed version
                         */
                        else
                        {
                            inst.gip_ins_class = gip_ins_class_store;
                            inst.gip_ins_subclass = ldm_stm_gip_ins_subclass;
                            inst.a = 1;
                            inst.s_or_stack = (alu_rn==13);
                            inst.p_or_offset_is_shift = 0;

                            inst.gip_ins_rm = arm_mapped_bottom_bit_set;
                            inst.gip_ins_rd = {type=gip_ins_r_type_none};
                            inst.gip_ins_rn = arm_mapped_rn;
                            inst.k = ldm_stm_num_regs[4;0]-1;

                            inst.valid = 1;

                            if (ldm_stm_num_regs==1)
                            {
                                next_cycle_of_opcode = 0;
                                pc_op = gip_pc_op_sequential;
                                if (ld_st_wb)
                                {
                                    inst.gip_ins_rd = arm_mapped_rn;
                                }
                            }
                            else
                            {
                                next_cycle_of_opcode[5;0] = ldm_stm_num_regs-2;
                                next_cycle_of_opcode[4] = 1;
                                pc_op = gip_pc_op_hold;
                            }

                            next_stored_reg_set[ldm_stm_bottom_bit_set] = 0;

                        }
                    }
                    /*b Handle later cycles - generate a 'ISTRCPA[S][F] #i (Acc), #+4 [->Rn] or preindexed version
                     */
                    else
                    {
                        inst.gip_ins_class = gip_ins_class_store;
                        inst.gip_ins_subclass = ldm_stm_gip_ins_subclass;
                        inst.gip_ins_cc = gip_ins_cc_cp;
                        inst.a = 1;
                        inst.s_or_stack = (alu_rn==13);
                        inst.p_or_offset_is_shift = 0;

                        inst.gip_ins_rm = arm_mapped_bottom_bit_set;
                        inst.gip_ins_rd = {type=gip_ins_r_type_none};
                        inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_acc};
                        inst.k = cycle_of_opcode[4;0];

                        inst.valid = 1;

                        if (cycle_of_opcode[4;0]==0) // No more to do after this one
                        {
                            next_cycle_of_opcode = 0;
                            pc_op = gip_pc_op_sequential;
                            if (ld_st_wb && ld_st_up)
                            {
                                inst.gip_ins_rd = arm_mapped_rn;
                            }
                        }
                        else
                        {
                            next_cycle_of_opcode[4] = 1;
                            next_cycle_of_opcode[4;0] = cycle_of_opcode[4;0]-1;
                            pc_op = gip_pc_op_hold;
                        }

                        next_stored_reg_set[ldm_stm_bottom_bit_set] = 0;

                    }

                    /*b However, if there are no registers in the original list, just ditch everything
                     */
                    if (ldm_stm_num_regs==0)
                    {
                        inst.valid = 0;
                        next_cycle_of_opcode = 0;
                        pc_op = gip_pc_op_sequential;
                    }
                }
                /*b Multiply
                 */
                case arm_ins_class_mul:
                {
                    full_switch (cycle_of_opcode)
                        {
                        case 0: /*b First the INIT instruction
                                 */
                        {
                            inst.gip_ins_class = gip_ins_class_arith;
                            inst.gip_ins_subclass = gip_ins_subclass_arith_init;
                            inst.a = 1;
                            inst.s_or_stack = 0;
                            inst.p_or_offset_is_shift = 1; // P required for INIT instruction

                            inst.gip_ins_rd = {type=gip_ins_r_type_none};
                            inst.gip_ins_rn = arm_mapped_rm; // Note reversal of rn and rm, and rn comes from rd!
                            inst.gip_ins_rm = arm_mapped_rd; // Note reversal of rn and rm, and rn comes from rd!
                            inst.immediate = 0;
                            if (opcode[21]) // Accumulate
                            {
                                inst.rm_is_imm = 0;
                            }
                            else
                            {
                                inst.rm_is_imm = 1;
                            }

                            inst.valid = 1;

                            next_cycle_of_opcode = 31;
                            pc_op = gip_pc_op_hold;
                        }
                        case 31: /*b Then the MLA instruction to get the ALU inputs ready, and do the first step
                                  */
                        {
                            inst.gip_ins_class = gip_ins_class_arith;
                            inst.gip_ins_subclass = gip_ins_subclass_arith_mla;
                            inst.gip_ins_cc = gip_ins_cc_cp;
                            inst.a = 1;
                            inst.s_or_stack = 0;
                            inst.p_or_offset_is_shift = 1; // P required for MLA instruction

                            inst.gip_ins_rd = {type=gip_ins_r_type_none};
                            inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_acc};
                            inst.gip_ins_rm = arm_mapped_rs;
                            inst.rm_is_imm = 0;

                            inst.valid = 1;

                            next_cycle_of_opcode = 30;
                            pc_op = gip_pc_op_hold;
                        }
                        case 30: /*b Then 14 MLB instruction to churn
                                  */
                        case 29:
                        case 28:
                        case 27:
                        case 26:
                        case 25:
                        case 24:
                        case 23:
                        case 22:
                        case 21:
                        case 20:
                        case 19:
                        case 18:
                        case 17:
                        {
                            inst.gip_ins_class = gip_ins_class_arith;
                            inst.gip_ins_subclass = gip_ins_subclass_arith_mlb;
                            inst.gip_ins_cc = gip_ins_cc_cp;
                            inst.a = 1;
                            inst.s_or_stack = 0;
                            inst.p_or_offset_is_shift = 1; // P required for MLA instruction

                            inst.gip_ins_rd = {type=gip_ins_r_type_none};
                            inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_acc};
                            inst.gip_ins_rm = arm_mapped_rs;
                            inst.immediate = 0;
                            inst.rm_is_imm = 1;

                            inst.valid = 1;

                            next_cycle_of_opcode = cycle_of_opcode-1;
                            pc_op = gip_pc_op_hold;
                        }
                        case 16: /*b Then the last MLB instruction to write the result
                                  */
                        {
                            inst.gip_ins_class = gip_ins_class_arith;
                            inst.gip_ins_subclass = gip_ins_subclass_arith_mlb;
                            inst.gip_ins_cc = gip_ins_cc_cp;
                            inst.a = 1;
                            inst.s_or_stack = 0;
                            inst.p_or_offset_is_shift = 1; // P required (?) for MLB instruction

                            inst.gip_ins_rd = arm_mapped_rn; // Note that rn contains rn... weird
                            inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_acc};
                            inst.gip_ins_rm = arm_mapped_rs;
                            inst.immediate = 0;
                            inst.rm_is_imm = 1;

                            inst.valid = 1;

                            next_cycle_of_opcode = 0;
                            pc_op = gip_pc_op_sequential;
                        }
                        }

                }
                /*b Branch
                 */
                case arm_ins_class_branch:
                {
                    /*b Handle 5 cases; conditional or not, link or not; split conditional branches to predicted or not, also
                     */
                    if (!branch_link)
                    {
                        if (!conditional) // guaranteed branch
                        {
                            inst.valid = 0;
                            pc_op = gip_pc_op_branch;
                            next_cycle_of_opcode = 0;
                        }
                        else
                        {
                            if (opcode[23]) // backward conditional branch; sub(!cc)f pc, #4 -> pc
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = gip_ins_subclass_arith_sub;
                                inst.gip_ins_cc = inv_cc;
                                inst.a = 0;
                                inst.s_or_stack = 0;
                                inst.p_or_offset_is_shift = 0;
                                inst.f = 1;
                                inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc};
                                inst.gip_ins_rd = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc};
                                inst.rm_is_imm = 1;
                                inst.immediate = 4;

                                inst.valid = 1;

                                pc_op = gip_pc_op_branch;
                                next_cycle_of_opcode = 0;
                            }
                            else // forward conditional branch; add[cc]f pc, #branch_offset -> pc
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = gip_ins_subclass_arith_add;
                                inst.a = 0;
                                inst.s_or_stack = 0;
                                inst.p_or_offset_is_shift = 0;
                                inst.f = 1;
                                inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc};
                                inst.gip_ins_rd = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc};
                                inst.rm_is_imm = 1;
                                inst.immediate = arm_branch_offset;

                                inst.valid = 1;

                                pc_op = gip_pc_op_sequential;
                                next_cycle_of_opcode = 0;
                            }
                        }
                    }
                    else
                    {
                        if (!conditional) // guaranteed branch with link; sub pc, #4 -> r14
                        {
                            inst.gip_ins_class = gip_ins_class_arith;
                            inst.gip_ins_subclass = gip_ins_subclass_arith_sub;
                            inst.a = 0;
                            inst.s_or_stack = 0;
                            inst.p_or_offset_is_shift = 0;
                            inst.f = 0;
                            inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc};
                            inst.gip_ins_rd = {type=gip_ins_r_type_register, r=14}; // Should map this
                            inst.rm_is_imm = 1;
                            inst.immediate = 4;

                            inst.valid = 1;

                            pc_op = gip_pc_op_branch;
                            next_cycle_of_opcode = 0;
                        }
                        else // conditional branch with link; sub{!cc}f pc, #4 -> pc; sub pc, #4 -> r14
                        {
                            full_switch (cycle_of_opcode)
                            {
                            case 0:
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = gip_ins_subclass_arith_sub;
                                inst.gip_ins_cc = inv_cc;
                                inst.a = 0;
                                inst.s_or_stack = 0;
                                inst.p_or_offset_is_shift = 0;
                                inst.f = 1;
                                inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc};
                                inst.gip_ins_rd = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc};
                                inst.rm_is_imm = 1;
                                inst.immediate = 4;

                                inst.valid = 1;

                                pc_op = gip_pc_op_hold;
                                next_cycle_of_opcode = 1;
                            }
                            default:
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = gip_ins_subclass_arith_sub;
                                inst.a = 0;
                                inst.s_or_stack = 0;
                                inst.p_or_offset_is_shift = 0;
                                inst.f = 0;
                                inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc};
                                inst.gip_ins_rd = {type=gip_ins_r_type_register, r=14}; // Should map this
                                inst.rm_is_imm = 1;
                                inst.immediate = 4;

                                inst.valid = 1;

                                pc_op = gip_pc_op_branch;
                                next_cycle_of_opcode = 0;
                            }
                            }
                        }
                    }

                }
                /*b Native
                 */
                case arm_ins_class_native:
                {
                    inst.gip_ins_cc = ins_cc;
                    next_cycle_of_opcode = 0;
                    pc_op = gip_pc_op_sequential;
                    arm_use_native_decode = 1;
                }
                /*b Done all instructions
                 */
                }

            /*b If condition is 'never' then just invalidate and ask for sequential!
             */
            if (cc==4hf)
            {
                inst.valid = 0;
                next_cycle_of_opcode = 0;
                pc_op = gip_pc_op_sequential;
            }

        }

    /*b Done
     */
}
