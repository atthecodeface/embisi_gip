/*a Copyright Gavin J Stark, 2004
 */

/*a To do
 */

/*a Constants
 */
constant integer max_requests = 4;
constant integer log_max_requests = 2;

/*a Types
 */

/*a fifo_ctrl_arb
 */
module fifo_ctrl_arb( input bit[max_requests] requests_in "Requests in",
                      output bit[max_requests] acknowledge_out "Acknowledges out; one will be asserted if at least one request is asserted; these are purely combinatorial",
                      output bit[log_max_requests] grant_to "Grant indicating which request is granted",
                      output bit granted "Asserted to indicate that a request is being handled" )

    /*b Documentation
     */
    "
This module implements a simple priority encoder to arbitrate between requesters for the FIFO

"
{

    /*b Aribter code
     */
    arbiter "Arbiter code":
        {
            acknowledge_out = 0;
            granted = 0;
            grant_to = 0;
            for ( i; max_requests )
            {
                if (requests_in[i])
                {
                    grant_to = i;
                    granted = 1;
                }
            }
            if (granted)
            {
                acknowledge_out[grant_to] = 1;
            }
        }
}
