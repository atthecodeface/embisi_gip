/*a Includes
 */
include "gip.h"
include "gip_internal.h"

/*a Types
 */

