/*a Includes
 */
include "gip.h"

/*a Module
 */
module gip_special( clock gip_clock,
                    input bit gip_reset,

                    input bit read,
                    input bit flush,
                    input bit[5] read_address,
                    output bit[32] read_data,
                    input bit write,
                    input bit[5] write_address,
                    input bit[32] write_data,

                    input bit[3] sched_state_thread,
                    input bit[4] sched_thread_data_config,
                    input bit[4] sched_thread_data_flag_dependencies,
                    input bit[32] sched_thread_data_pc,

                    input bit[5] postbus_semaphore_to_set "Semaphore to set due to postbus receive/transmit - none if zero",

                    output bit[8] special_repeat_count,
                    output bit[2] special_alu_mode,
                    output bit special_cp_trail_2,
                    output bit[32] special_semaphores,
                    output bit special_cooperative,
                    output bit special_round_robin,
                    output bit special_thread_data_write_pc,
                    output bit special_thread_data_write_config,
                    output bit[3] special_write_thread,
                    output bit[32] special_thread_data_pc,
                    output bit[4] special_thread_data_config,
                    output bit[4] special_thread_data_flag_dependencies,
                    output bit[3] special_selected_thread

    )
{
    /*b Default clock and reset
     */
    default clock gip_clock;
    default reset gip_reset;

    /*b State in the special registers guaranteed by the design
     */
    clocked bit[32] special_semaphores = 1;
    clocked bit[32] special_semaphores_mask = 0; // semaphores to set/clear on next sempahore read
    clocked bit special_cooperative = 0;
    clocked bit special_round_robin = 0;
    clocked bit thread_0_privilege = 0;
    clocked bit[3] special_selected_thread = 0; // Thread to read or write
    clocked bit[3] special_write_thread = 0; // Thread to actually use for writing thread_data_pc/config
    clocked bit special_thread_data_write_pc = 0; // 1 if the thread_data_pc should be written to write_thread
    clocked bit special_thread_data_write_config = 0; // 1 if the thread_data_config should be written to write_thread
    clocked bit[32] special_thread_data_pc = 0;
    clocked bit[4] special_thread_data_config = 0;
    clocked bit[4] special_thread_data_flag_dependencies = 0;
    clocked bit[8] special_repeat_count=0; // repeat count
    clocked bit[5] arm_trap_semaphore = 0;

    clocked bit[32] preempted_pc_l=0;
    clocked bit[32] preempted_pc_m=0;
    clocked bit[4] preempted_flags_l=0;
    clocked bit[4] preempted_flags_m=0;

    /*b Combinatorials
     */
    comb bit[32]new_semaphores;

    /*b NYI
     */
    nyi "":
        {
            special_cp_trail_2 = special_repeat_count[0];
            special_alu_mode = special_repeat_count[2;0];
        }
    /*b Read process
     */
    read_process "Read the special registers":
    {
        read_data = 0;
        if (read)
        {
            part_switch (read_address)
                {
                case gip_special_reg_semaphores_set:
                case gip_special_reg_semaphores_clear:
                {
                    read_data = special_semaphores;
                }
                case gip_special_reg_thread:
                {
                    read_data[3;0] = special_selected_thread;
                }
                case gip_special_reg_thread_pc:
                {
                    read_data = special_thread_data_pc;
                }
                case gip_special_reg_thread_data:
                {
                    read_data[4;0] = special_thread_data_config;
                    read_data[4;4] = special_thread_data_flag_dependencies;
                }
                case gip_special_reg_preempted_pc_l:
                {
                    read_data = preempted_pc_l;
                }
                case gip_special_reg_preempted_pc_m:
                {
                    read_data = preempted_pc_l;
                }
                case gip_special_reg_preempted_flags_l:
                {
                    read_data[4;0] = preempted_flags_l;
                }
                case gip_special_reg_preempted_flags_m:
                {
                    read_data[4;0] = preempted_flags_m;
                }
                }
        }
    }

    /*b Write process
     */
    write_process "Write the special registers":
    {
        /*b Default values for interacting with scheduler
         */
        special_thread_data_write_pc <= 0;
        special_thread_data_write_config <= 0;
        special_thread_data_pc <= sched_thread_data_pc;
        special_thread_data_config <= sched_thread_data_config;
        special_thread_data_flag_dependencies <= sched_thread_data_flag_dependencies;
        special_write_thread <= special_selected_thread;

        /*b Handle writes
         */
        if (write)
        {
            part_switch (write_address)
                {
                case gip_special_reg_gip_config:
                {
                    special_cooperative <= write_data[0];
                    special_round_robin <= write_data[1];
                    thread_0_privilege <= write_data[2];
                    arm_trap_semaphore <= write_data[5;16];
                }
                case gip_special_reg_semaphores_set:
                case gip_special_reg_semaphores_clear:
                {
                    special_semaphores_mask <= write_data;
                }
                case gip_special_reg_thread:
                {
                    special_selected_thread <= write_data[3;0];
                }
                case gip_special_reg_thread_pc:
                {
                    special_thread_data_write_pc <= 1;
                    special_thread_data_pc[0] <= 0;
                    special_thread_data_pc[31;1] <= write_data[31;1];
                    if (write_data[0])
                    {
                        special_write_thread <= special_selected_thread;
                    }
                    else
                    {
                        special_write_thread <= sched_state_thread;
                    }
                }
                case gip_special_reg_thread_data:
                {
                    special_thread_data_write_config <= 1;
                    special_thread_data_config <= write_data[4;0];
                    special_thread_data_flag_dependencies <= write_data[4;4];
                    if (write_data[8])
                    {
                        special_write_thread <= special_selected_thread;
                    }
                    else
                    {
                        special_write_thread <= sched_state_thread;
                    }
                }
                case gip_special_reg_repeat_count:
                {
                    special_repeat_count <= write_data[8;0];
                }
                case gip_special_reg_preempted_pc_l:
                {
                    preempted_pc_l <= write_data;
                }
                case gip_special_reg_preempted_pc_m:
                {
                    preempted_pc_m <= write_data;
                }
                case gip_special_reg_preempted_flags_l:
                {
                    preempted_flags_l <= write_data[4;0];
                }
                case gip_special_reg_preempted_flags_m:
                {
                    preempted_flags_m <= write_data[4;0];
                }
                }
        }

        /*b Handle setting and clearing of semaphores
         */
        new_semaphores = special_semaphores;
        if (read && !flush)
        {
            if (read_address==gip_special_reg_semaphores_clear)
            {
                special_semaphores_mask <= 0;
                new_semaphores = special_semaphores &~ special_semaphores_mask;
            }
            if (read_address==gip_special_reg_semaphores_set)
            {
                special_semaphores_mask <= 0;
                new_semaphores = special_semaphores | special_semaphores_mask;
            }
        }
        if (postbus_semaphore_to_set)
        {
            new_semaphores[postbus_semaphore_to_set] = 1;
        }

        /*b Set semaphores
         */
        special_semaphores <= new_semaphores;
    }

    /*b Done
     */
}

