/*a Copyright Gavin J Stark, 2004
 */

/*a To do
 */

/*a Constants
 */
constant integer max_requests = 4;
constant integer log_max_requests = 2;

/*a Types
 */

/*a fifo_ctrl_arb
 */
module fifo_ctrl_arb( input bit[max_requests] requests_in "Requests in",
                      output bit[max_requests] acknowledge_out "Acknowledges out; one will be asserted if at least one request is asserted; these are purely combinatorial",
                      output bit[log_max_requests] grant_to "Grant indicating which request is granted",
                      output bit granted "Asserted to indicate that a request is being handled" )

    /*b Documentation
     */
    "
This module implements a simple priority encoder to arbitrate between requesters for the FIFO

"
{

    /*b Aribter code
     */
    arbiter "Arbiter code":
        {
            acknowledge_out = 0;
            granted = 0;
            grant_to = 0;
            if (requests_in[0])
            {
                acknowledge_out[0] = 1;
                grant_to = 0;
                granted = 1;
            }
            elsif (requests_in[1])
                {
                    acknowledge_out[1] = 1;
                    grant_to = 1;
                    granted = 1;
                }
            elsif (requests_in[2])
                {
                    acknowledge_out[2] = 1;
                    grant_to = 2;
                    granted = 1;
                }
            elsif (requests_in[3])
                {
                    acknowledge_out[3] = 1;
                    grant_to = 3;
                    granted = 1;
                }
        }
}
