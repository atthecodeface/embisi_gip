/*a Includes
 */
include "gip.h"
include "gip_internal.h"

/*a Types
 */

/*a Module
 */
module gip_decode_native( input bit[16] opcode,

                          input bit[8] special_repeat_count,
                          input bit[2] special_alu_mode,

                          output t_gip_instruction_rf inst,
                          output t_gip_pc_op pc_op,
                          output bit[32] native_mapped_branch_offset,

                          input bit extended,
                          input bit[28] extended_immediate,
                          input t_gip_ins_r extended_rd,
                          input t_gip_ins_r extended_rn,
                          input t_gip_ins_r extended_rm,
                          input t_gip_ext_cmd extended_cmd,

                          output bit extending,
                          output bit[28] next_extended_immediate,
                          output t_gip_ins_r next_extended_rd,
                          output t_gip_ins_r next_extended_rn,
                          output t_gip_ins_r next_extended_rm,
                          output t_gip_ext_cmd next_extended_cmd,

                          output bit[6] next_atomic,

                          input bit in_conditional_shadow,
                          input bit in_immediate_conditional_shadow,
                          output bit next_in_immediate_conditional_shadow

                          )
{
    comb bit[4] ins_class;
    comb bit[4] ins_subclass;
    comb bit[5] ins_subclass_full;
    comb bit[3] ins_subclass_ldst;
    comb bit[2] ins_subclass_shift;
    comb bit[8] full_rd;
    comb bit[4] rd;
    comb bit[4] rn;
    comb bit[4] rm;
    comb bit[4] imm;
    comb bit[4] cond;
    comb bit sign;
    comb bit acc;
    comb bit[2] op;
    comb bit[4] burst;
    comb bit shift_is_imm;
    comb bit[5] shift_imm;
    comb bit branch_delay_slot;
    comb bit[32] branch_offset;
    comb bit store_not_load;

    comb t_gip_ins_r native_mapped_rd;
    comb bit native_mapped_rd_is_pc;
    comb t_gip_ins_r native_mapped_rn;
    comb t_gip_ins_r native_mapped_rm;
    comb t_gip_ins_r native_mapped_rm_full_extend;
    comb bit[32] native_mapped_immediate;

    comb bit[2] alu_mode;

    /*b Break out instruction
     */
    breakout_instruction "Breakout instruction":
        {
            ins_class = opcode[4;12]; // instruction class
            ins_subclass = opcode[4;8]; // instruction subclass for ALU, cond instructions
            ins_subclass_shift = opcode[2;10]; // instruction subclass for shift instructions
            full_rd = opcode[8;4]; // full extension of rd for ext instructions
            rm = opcode[4;0]; // rm for nonextended instructions (ALU, cond) and extrnm, extrdrm; data register for loads and stores
            rd = opcode[4;4]; // rd for nonextended instructions (ALU, cond); address for loads and stores
            rn = opcode[4;8]; // rn for extrnm (nonextended instructions are 2-register)
            imm = opcode[4;0];// 4 bit immediate for not extimm instructions (ALU, cond)
            cond = opcode[4;8]; // 4 bit cond for extcmd
            sign = opcode[7]; // 1 bit sign for extcmd
            acc = opcode[6]; // 1 bit acc for extcmd
            op = opcode[2;4]; // 2 bit options for extcmd
            burst = opcode[4;0]; // 4 bit burst for extcmd

            shift_is_imm = opcode[9];
            shift_imm[4;0] = opcode[4;0];
            shift_imm[4] = opcode[8];

            branch_delay_slot = opcode[0];
            branch_offset = 0;
            branch_offset[11;1] = opcode[11;1];
            if (opcode[11])
            {
                branch_offset[20;12] = -1;
            }

            store_not_load = opcode[8];
            ins_subclass_ldst = opcode[3;9];
        }

    /*b Map registers and immediate
     */
    map_registers "Map registers and immediate value using the extended amounts in the current registers (from previous instruction decodes)":
        {
            /*b Map rd to instruction rd; pc if that is 15; but if extended, to full given extension
             */
            native_mapped_rd.type = gip_ins_r_type_register;
            native_mapped_rd.r = 0;
            native_mapped_rd.r[4;0] = rd;
            if (rd==15) { native_mapped_rd = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc}; }
            if (extended_rd.type!=gip_ins_r_type_no_override) { native_mapped_rd = extended_rd; }
            native_mapped_rd_is_pc = ( (native_mapped_rd.type==gip_ins_r_type_internal) &&
                                       (native_mapped_rd.r==gip_ins_r_int_pc) );

            /*b Map rn to instruction rd; acc if that is 15; but if extended, to full given extension
             */
            native_mapped_rn.type = gip_ins_r_type_register;
            native_mapped_rn.r = 0;
            native_mapped_rn.r[4;0] = rd;
            if (rd==15) { native_mapped_rn = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_acc}; }
            if (extended_rn.type!=gip_ins_r_type_no_override) { native_mapped_rn = extended_rn; }

            /*b Map rm to instruction rm; pc if that is 15; but if extended, to full given extension
             */
            native_mapped_rm.type = gip_ins_r_type_register;
            native_mapped_rm.r = 0;
            native_mapped_rm.r[4;0] = rm;
            if (rm==15) { native_mapped_rm = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_acc}; }
            native_mapped_rm_full_extend = native_mapped_rm;
            if (extended_rm.type!=gip_ins_r_type_no_override)
            {
                native_mapped_rm_full_extend = extended_rm;
                native_mapped_rm.type = extended_rm.type;
                native_mapped_rm.r[4]=extended_rm.r[4];
                native_mapped_rm.r[4;0]=rm;
            }

            /*b Map the immediate value in the instruction
             */
            native_mapped_immediate[28;4] = extended_immediate;
            native_mapped_immediate[4;0] = imm;

            /*b Map the branch offset
             */
            native_mapped_branch_offset = branch_offset;
            if (extended_immediate!=0)
            {
                native_mapped_branch_offset[20;12] = extended_immediate[20;0];
            }
            native_mapped_branch_offset[12;0] = branch_offset[12;0];
        }

    /*b Decode instruction
     */
    decode_instruction "Decode instruction":
        {
            /*b Define outputs as a NOP
             */
            pc_op = gip_pc_op_sequential;
            next_extended_immediate = extended_immediate;
            next_extended_rd = {type=gip_ins_r_type_no_override, r=0};
            next_extended_rm = {type=gip_ins_r_type_no_override, r=0};
            next_extended_rn = {type=gip_ins_r_type_no_override, r=0};
            next_extended_cmd = {extended=0, cc=gip_ins_cc_always, sign_or_stack=0, acc=0, op=0, burst=0};
            extending = 0;
            next_in_immediate_conditional_shadow = 0;
            next_atomic = 0;

            inst.gip_ins_class = gip_ins_class_logic;
            inst.gip_ins_subclass = gip_ins_subclass_logic_mov;
            inst.gip_ins_cc = gip_ins_cc_always;
            inst.a = 0;
            inst.s_or_stack = 0;
            inst.p_or_offset_is_shift = 0;
            inst.k = 0;
            inst.f = 0;
            inst.d = 0;
            inst.gip_ins_rm = native_mapped_rm;
            inst.gip_ins_rn = native_mapped_rn;
            inst.rm_is_imm = 0;
            inst.immediate = native_mapped_immediate;
            inst.gip_ins_rd = native_mapped_rd;
            inst.tag = 0;
            inst.valid = 0;

            if (extended_cmd.extended)
            {
                inst.a = extended_cmd.acc;
                inst.s_or_stack = extended_cmd.sign_or_stack;
                if (extended_cmd.cc!=14)
                {
                    inst.gip_ins_cc = extended_cmd.cc;
                }
            }

            /*b Decode instruction according to class
             */
            full_switch (ins_class)
                {
                /*b Debug
                 */
                case gip_native_ins_class_debug: // Debug - do nothing for now
                {
                    pc_op = gip_pc_op_sequential;
                }
                /*b Extimm (4)
                 */
                case gip_native_ins_class_extimm_0:
                case gip_native_ins_class_extimm_1:
                case gip_native_ins_class_extimm_2:
                case gip_native_ins_class_extimm_3:
                {
                    if (extended_immediate==0)
                    {
                        next_extended_immediate[14;0] = opcode[14;0];
                        if (opcode[13])
                        {
                            next_extended_immediate[14;14] = -1;
                        }
                    }
                    else
                    {
                        next_extended_immediate[14;14] = extended_immediate[14;0];
                        next_extended_immediate[14;0] = opcode[14;0];
                    }
                    extending = 1;
                }
                /*b Extrdrm
                 */
                case gip_native_ins_class_extrdrm:
                {
                    next_extended_rd.type = full_rd[3;5];
                    next_extended_rd.r = full_rd[5;0];
                    next_extended_rm.type = rm[3;1];
                    next_extended_rm.r = 0;
                    next_extended_rm.r[4] = rm[0];
                    extending = 1;
                }
                /*b Extrnrm
                 */
                case gip_native_ins_class_extrnrm:
                {
                    next_extended_rn.type = rn[3;1];
                    next_extended_rn.r = 0;
                    next_extended_rn.r[4] = rn[0];
                    next_extended_rm.type = rm[3;1];
                    next_extended_rm.r = 0;
                    next_extended_rm.r[4] = rm[0];
                    extending = 1;
                }
                /*b Extcmd
                 */
                case gip_native_ins_class_extcmd:
                {
                    next_extended_cmd.extended = 1;
                    next_extended_cmd.cc = cond;
                    next_extended_cmd.sign_or_stack = sign;
                    next_extended_cmd.acc = acc;
                    next_extended_cmd.op = op;
                    next_extended_cmd.burst = burst;
                }
                /*b ALU (reg and imm)
                 */
                case gip_native_ins_class_alu_reg:
                case gip_native_ins_class_alu_imm:
                {
                    /*b Decode mode and ALU operations
                     */
                    alu_mode = special_alu_mode;
                    if (extended_cmd.extended)
                    {
                        if (extended_cmd.op!=0)
                        {
                            alu_mode = extended_cmd.op;
                        }
                    }
                    else
                    {
                        inst.a = 1;
                        inst.s_or_stack = 1;
                    }
                    /*b Basic instructions - get inst.gip_ins_class and inst.gip_ins_subclass
                     */
                    if (!ins_subclass[3])
                    {
                        part_switch (ins_subclass)
                        {
                        case gip_native_ins_subclass_alu_and:
                        {
                            inst.gip_ins_class = gip_ins_class_logic;
                            inst.gip_ins_subclass = gip_ins_subclass_logic_and;
                        }
                        case gip_native_ins_subclass_alu_or:
                        {
                            inst.gip_ins_class = gip_ins_class_logic;
                            inst.gip_ins_subclass = gip_ins_subclass_logic_or;
                        }
                        case gip_native_ins_subclass_alu_xor:
                        {
                            inst.gip_ins_class = gip_ins_class_logic;
                            inst.gip_ins_subclass = gip_ins_subclass_logic_xor;
                        }
                        case gip_native_ins_subclass_alu_mov:
                        {
                            inst.gip_ins_class = gip_ins_class_logic;
                            inst.gip_ins_subclass = gip_ins_subclass_logic_mov;
                        }
                        case gip_native_ins_subclass_alu_mvn:
                        {
                            inst.gip_ins_class = gip_ins_class_logic;
                            inst.gip_ins_subclass = gip_ins_subclass_logic_mvn;
                        }
                        case gip_native_ins_subclass_alu_add:
                        {
                            inst.gip_ins_class = gip_ins_class_arith;
                            inst.gip_ins_subclass = gip_ins_subclass_arith_add;
                        }
                        case gip_native_ins_subclass_alu_sub:
                        {
                            inst.gip_ins_class = gip_ins_class_arith;
                            inst.gip_ins_subclass = gip_ins_subclass_arith_sub;
                        }
                        case gip_native_ins_subclass_alu_adc:
                        {
                            inst.gip_ins_class = gip_ins_class_arith;
                            inst.gip_ins_subclass = gip_ins_subclass_arith_adc;
                        }
                        }
                    }
                    /*b Modal instructions
                     */
                    else
                    {
                        part_switch (alu_mode)
                        {
                            /*b Bit mode
                             */
                        case gip_native_mode_bit:
                        {
                            part_switch (ins_subclass)
                            {
                            case gip_native_ins_subclass_alu_xorfirst:
                            {
                                inst.gip_ins_class = gip_ins_class_logic;
                                inst.gip_ins_subclass = gip_ins_subclass_logic_xorfirst;
                            }
                            case gip_native_ins_subclass_alu_rsb:
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = gip_ins_subclass_arith_rsb;
                            }
                            case gip_native_ins_subclass_alu_bic:
                            {
                                inst.gip_ins_class = gip_ins_class_logic;
                                inst.gip_ins_subclass = gip_ins_subclass_logic_bic;
                            }
                            case gip_native_ins_subclass_alu_orn:
                            {
                                inst.gip_ins_class = gip_ins_class_logic;
                                inst.gip_ins_subclass = gip_ins_subclass_logic_orn;
                            }
                            case gip_native_ins_subclass_alu_andcnt:
                            {
                                inst.gip_ins_class = gip_ins_class_logic;
                                inst.gip_ins_subclass = gip_ins_subclass_logic_andcnt;
                            }
                            case gip_native_ins_subclass_alu_xorlast:
                            {
                                inst.gip_ins_class = gip_ins_class_logic;
                                inst.gip_ins_subclass = gip_ins_subclass_logic_xorlast;
                            }
                            case gip_native_ins_subclass_alu_bitreverse:
                            {
                                inst.gip_ins_class = gip_ins_class_logic;
                                inst.gip_ins_subclass = gip_ins_subclass_logic_bitreverse;
                            }
                            case gip_native_ins_subclass_alu_bytereverse:
                            {
                                inst.gip_ins_class = gip_ins_class_logic;
                                inst.gip_ins_subclass = gip_ins_subclass_logic_bytereverse;
                            }
                            }
                        }
                            /*b Math mode
                             */
                        case gip_native_mode_math:
                        {
                            part_switch (ins_subclass)
                            {
                            case gip_native_ins_subclass_alu_xorfirst:
                            {
                                inst.gip_ins_class = gip_ins_class_logic;
                                inst.gip_ins_subclass = gip_ins_subclass_logic_xorfirst;
                            }
                            case gip_native_ins_subclass_alu_rsb:
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = gip_ins_subclass_arith_rsb;
                            }
                            case gip_native_ins_subclass_alu_init:
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = gip_ins_subclass_arith_init;
                            }
                            case gip_native_ins_subclass_alu_mla:
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = gip_ins_subclass_arith_mla;
                            }
                            case gip_native_ins_subclass_alu_mlb:
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = gip_ins_subclass_arith_mlb;
                            }
                            case gip_native_ins_subclass_alu_sbc:
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = gip_ins_subclass_arith_sbc;
                            }
                            case gip_native_ins_subclass_alu_dva:
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = gip_ins_subclass_arith_dva;
                            }
                            case gip_native_ins_subclass_alu_dvb:
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = gip_ins_subclass_arith_dvb;
                            }
                            }
                        }
                            /*b GP mode
                             */
                        case gip_native_mode_gp:
                        {
                            part_switch (ins_subclass)
                            {
                            case gip_native_ins_subclass_alu_xorfirst:
                            {
                                inst.gip_ins_class = gip_ins_class_logic;
                                inst.gip_ins_subclass = gip_ins_subclass_logic_xorfirst;
                            }
                            case gip_native_ins_subclass_alu_rsb:
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = gip_ins_subclass_arith_rsb;
                            }
                            case gip_native_ins_subclass_alu_bic:
                            {
                                inst.gip_ins_class = gip_ins_class_logic;
                                inst.gip_ins_subclass = gip_ins_subclass_logic_bic;
                            }
                            case gip_native_ins_subclass_alu_andxor:
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = gip_ins_subclass_logic_andxor;
                            }
                            case gip_native_ins_subclass_alu_rsc:
                            {
                                inst.gip_ins_class = gip_ins_class_arith;
                                inst.gip_ins_subclass = gip_ins_subclass_arith_rsc;
                            }
                            }
                        }
                        }
                    }
                    /*b Map remains of instruction
                     */
                    inst.f = native_mapped_rd_is_pc;
                    if (ins_class==gip_native_ins_class_alu_imm)
                    {
                        inst.rm_is_imm = 1;
                        inst.gip_ins_rm.type = gip_ins_r_type_none;
                    }
                    else
                    {
                        inst.rm_is_imm = 0;
                    }
                    inst.valid = 1;
                }
                /*b Conditional instructions (reg and imm) 
                 */
                case gip_native_ins_class_cond_reg:
                case gip_native_ins_class_cond_imm:
                {
                    /*b Decode mode and operation, rd
                     */
                    ins_subclass_full = 0;
                    ins_subclass_full[4;0] = ins_subclass;
                    if (extended_cmd.extended)
                    {
                        ins_subclass_full[4] = extended_cmd.op[0]; // use op bit 0 as top bit of conditional
                    }
                    else
                    {
                        inst.a = 1;
                        inst.s_or_stack = 0;
                        inst.gip_ins_cc = gip_ins_cc_always; // Unless in AND mode and in direct shadow of a conditional, when it should be CP
                        if (in_immediate_conditional_shadow)
                        {
                            inst.gip_ins_cc = gip_ins_cc_cp;
                        }
                    }
                    /*b Get arithmetic operation for requested subclass
                     */
                    inst.gip_ins_class = gip_ins_class_arith;
                    inst.gip_ins_subclass = gip_ins_subclass_arith_sub;
                    part_switch (ins_subclass_full)
                        {
                        case gip_native_ins_subclass_cond_eq:
                        case gip_native_ins_subclass_cond_ne:
                        case gip_native_ins_subclass_cond_gt:
                        case gip_native_ins_subclass_cond_ge:
                        case gip_native_ins_subclass_cond_lt:
                        case gip_native_ins_subclass_cond_le:
                        case gip_native_ins_subclass_cond_hi:
                        case gip_native_ins_subclass_cond_hs:
                        case gip_native_ins_subclass_cond_lo:
                        case gip_native_ins_subclass_cond_ls:
                        case gip_native_ins_subclass_cond_seq:
                        case gip_native_ins_subclass_cond_sne:
                        case gip_native_ins_subclass_cond_sgt:
                        case gip_native_ins_subclass_cond_sge:
                        case gip_native_ins_subclass_cond_slt:
                        case gip_native_ins_subclass_cond_sle:
                        case gip_native_ins_subclass_cond_shi:
                        case gip_native_ins_subclass_cond_shs:
                        case gip_native_ins_subclass_cond_slo:
                        case gip_native_ins_subclass_cond_sls:
                        case gip_native_ins_subclass_cond_smi:
                        case gip_native_ins_subclass_cond_spl:
                        case gip_native_ins_subclass_cond_svs:
                        case gip_native_ins_subclass_cond_svc:
                        {
                            inst.gip_ins_class = gip_ins_class_arith;
                            inst.gip_ins_subclass = gip_ins_subclass_arith_sub;
                        }
                        case gip_native_ins_subclass_cond_sps:
                        case gip_native_ins_subclass_cond_spc:
                        {
                            inst.gip_ins_class = gip_ins_class_logic;
                            inst.gip_ins_subclass = gip_ins_subclass_logic_mov;
                            inst.p_or_offset_is_shift = 1;
                        }
                        case gip_native_ins_subclass_cond_allset:
                        case gip_native_ins_subclass_cond_anyclr:
                        {
                            inst.gip_ins_class = gip_ins_class_logic;
                            inst.gip_ins_subclass = gip_ins_subclass_logic_andxor;
                        }
                        case gip_native_ins_subclass_cond_allclr:
                        case gip_native_ins_subclass_cond_anyset:
                        {
                            inst.gip_ins_class = gip_ins_class_logic;
                            inst.gip_ins_subclass = gip_ins_subclass_logic_and;
                        }
                        }
                    /*b Get target condition
                     */
                    inst.gip_ins_rd.type = gip_ins_r_type_internal;
                    part_switch (ins_subclass_full)
                        {
                        case gip_native_ins_subclass_cond_eq:
                        case gip_native_ins_subclass_cond_allset:
                        case gip_native_ins_subclass_cond_allclr:
                        case gip_native_ins_subclass_cond_seq:
                        case gip_native_ins_subclass_cond_sne:
                        case gip_native_ins_subclass_cond_sgt:
                        case gip_native_ins_subclass_cond_sge:
                        case gip_native_ins_subclass_cond_slt:
                        case gip_native_ins_subclass_cond_sle:
                        case gip_native_ins_subclass_cond_shi:
                        case gip_native_ins_subclass_cond_shs:
                        case gip_native_ins_subclass_cond_slo:
                        case gip_native_ins_subclass_cond_sls:
                        case gip_native_ins_subclass_cond_smi:
                        case gip_native_ins_subclass_cond_spl:
                        case gip_native_ins_subclass_cond_svs:
                        case gip_native_ins_subclass_cond_svc:
                        {
                            inst.gip_ins_rd.r = gip_ins_rd_int_eq;
                        }
                        case gip_native_ins_subclass_cond_anyclr:
                        case gip_native_ins_subclass_cond_anyset:
                        case gip_native_ins_subclass_cond_ne:
                        {
                            inst.gip_ins_rd.r = gip_ins_rd_int_ne;
                        }
                        case gip_native_ins_subclass_cond_gt:
                        {
                            inst.gip_ins_rd.r = gip_ins_rd_int_gt;
                        }
                        case gip_native_ins_subclass_cond_ge:
                        {
                            inst.gip_ins_rd.r = gip_ins_rd_int_ge;
                        }
                        case gip_native_ins_subclass_cond_lt:
                        {
                            inst.gip_ins_rd.r = gip_ins_rd_int_lt;
                        }
                        case gip_native_ins_subclass_cond_le:
                        {
                            inst.gip_ins_rd.r = gip_ins_rd_int_le;
                        }
                        case gip_native_ins_subclass_cond_hi:
                        {
                            inst.gip_ins_rd.r = gip_ins_rd_int_hi;
                        }
                        case gip_native_ins_subclass_cond_hs:
                        case gip_native_ins_subclass_cond_sps:
                        {
                            inst.gip_ins_rd.r = gip_ins_rd_int_cs;
                        }
                        case gip_native_ins_subclass_cond_spc:
                        case gip_native_ins_subclass_cond_lo:
                        {
                            inst.gip_ins_rd.r = gip_ins_rd_int_cc;
                        }
                        case gip_native_ins_subclass_cond_ls:
                        {
                            inst.gip_ins_rd.r = gip_ins_rd_int_ls;
                        }
                        }
                    /*b Get conditional if override required
                     */
                    part_switch (ins_subclass_full)
                        {
                        case gip_native_ins_subclass_cond_seq:
                        {
                            inst.gip_ins_cc = gip_ins_cc_eq;
                        }
                        case gip_native_ins_subclass_cond_sne:
                        {
                            inst.gip_ins_cc = gip_ins_cc_ne;
                        }
                        case gip_native_ins_subclass_cond_sgt:
                        {
                            inst.gip_ins_cc = gip_ins_cc_gt;
                        }
                        case gip_native_ins_subclass_cond_sge:
                        {
                            inst.gip_ins_cc = gip_ins_cc_ge;
                        }
                        case gip_native_ins_subclass_cond_slt:
                        {
                            inst.gip_ins_cc = gip_ins_cc_lt;
                        }
                        case gip_native_ins_subclass_cond_sle:
                        {
                            inst.gip_ins_cc = gip_ins_cc_le;
                        }
                        case gip_native_ins_subclass_cond_shi:
                        {
                            inst.gip_ins_cc = gip_ins_cc_hi;
                        }
                        case gip_native_ins_subclass_cond_shs:
                        {
                            inst.gip_ins_cc = gip_ins_cc_cs;
                        }
                        case gip_native_ins_subclass_cond_slo:
                        {
                            inst.gip_ins_cc = gip_ins_cc_cc;
                        }
                        case gip_native_ins_subclass_cond_sls:
                        {
                            inst.gip_ins_cc = gip_ins_cc_ls;
                        }
                        case gip_native_ins_subclass_cond_smi:
                        {
                            inst.gip_ins_cc = gip_ins_cc_mi;
                        }
                        case gip_native_ins_subclass_cond_spl:
                        {
                            inst.gip_ins_cc = gip_ins_cc_pl;
                        }
                        case gip_native_ins_subclass_cond_svs:
                        {
                            inst.gip_ins_cc = gip_ins_cc_vs;
                        }
                        case gip_native_ins_subclass_cond_svc:
                        {
                            inst.gip_ins_cc = gip_ins_cc_vc;
                        }
                        }
                    /*b Map other
                     */
                    if (ins_class==gip_native_ins_class_cond_imm)
                    {
                        inst.rm_is_imm = 1;
                        inst.gip_ins_rm.type = gip_ins_r_type_none;
                    }
                    else
                    {
                        inst.rm_is_imm = 0;
                    }
                    inst.valid = 1;
                    next_in_immediate_conditional_shadow = 1;
                }
                /*b Shift instruction (subclasses lsr, asr, lsl, ror, with immediate/reg)
                 */
                case gip_native_ins_class_shift:
                {
                    /*b Decode shift operation
                     */
                    if (!extended_cmd.extended)
                    {
                        inst.s_or_stack = 1;
                    }
                    full_switch (ins_subclass_shift)
                    {
                    case gip_native_ins_subclass_shift_lsl:
                    {
                        inst.gip_ins_subclass = gip_ins_subclass_shift_lsl;
                    }
                    case gip_native_ins_subclass_shift_lsr:
                    {
                        inst.gip_ins_subclass = gip_ins_subclass_shift_lsr;
                    }
                    case gip_native_ins_subclass_shift_asr:
                    {
                        inst.gip_ins_subclass = gip_ins_subclass_shift_asr;
                    }
                    case gip_native_ins_subclass_shift_ror:
                    {
                        inst.gip_ins_subclass = gip_ins_subclass_shift_ror;
                        if (shift_is_imm && (shift_imm==0))
                        {
                            inst.gip_ins_subclass = gip_ins_subclass_shift_ror33;
                        }
                    }
                    }
                    inst.f = native_mapped_rd_is_pc;
                    if (shift_is_imm)
                    {
                        inst.rm_is_imm = 1;
                        inst.gip_ins_rm.type = gip_ins_r_type_none;
                    }
                    else
                    {
                        inst.rm_is_imm = 0;
                    }
                    inst.valid = 1;
                }
                /*b Memory instructions (subclasses are ldr and str)
                 */
                case gip_native_ins_class_memory:
                {
                    if (!store_not_load)
                    {
                        /*b Decode basic defaults for a load - ldr rd, address_mode(rn)
                         */
                        inst.rm_is_imm = 0;
                        // rm (offset to address to store) defaults to native_mapped_rm; we need the fully extended version if it is used as the instruction supplies no rm bits
                        // rn (address to store) defaults to native_mapped_rn
                        // rd (data to store) defaults to native_mapped_rd; this is only correct if native_mapped_rd picks up the (normally) 'rm' bits of the instruction opcode
                        // We actually have a choice here
                        //  data to read into could be native_mapped_rm
                        //       and offset could be extended rd
                        // or
                        //  data to read into could be native_mapped_rd, but change the source of rd bit in the instruction from 4;4 to 4;0
                        //       and offset could be native_mapped_rm_full_extend
                        // we actually use the former
                        // SO
                        //  gip_ins_rd = native_mapped_rm
                        //  gip_ins_rm = native_mapped_rd IF extended and if an index is required
                        if (!extended_cmd.extended)
                        {
                            inst.a = 1;
                            inst.s_or_stack = 0;
                        }
                        inst.k = 0;
                        inst.gip_ins_rd = native_mapped_rm; 
                        inst.gip_ins_rm = native_mapped_rd;
                        inst.gip_ins_class = gip_ins_class_load;
                        /*b Determine subclass for a load, and immediate value
                         */
                        full_switch (ins_subclass_ldst)
                        {
                        case gip_native_ins_subclass_memory_word_noindex: // Preindex Up Word, immediate of zero (unless extended - then preindex up by immediate value)
                        {
                            inst.gip_ins_subclass = gip_ins_subclass_memory_word | gip_ins_subclass_memory_up | gip_ins_subclass_memory_preindex;
                            inst.immediate[4;0] = 0;
                            inst.rm_is_imm = 1;
                            inst.gip_ins_rm.type = gip_ins_r_type_none;
                        }
                        case gip_native_ins_subclass_memory_half_noindex: // Preindex Up Half, immediate of zero (unless extended - then preindex up by immediate value)
                        {
                            inst.gip_ins_subclass = gip_ins_subclass_memory_half | gip_ins_subclass_memory_up | gip_ins_subclass_memory_preindex;
                            inst.immediate[4;0] = 0;
                            inst.rm_is_imm = 1;
                            inst.gip_ins_rm.type = gip_ins_r_type_none;
                        }
                        case gip_native_ins_subclass_memory_byte_noindex: // Preindex Up Byte, immediate of zero (unless extended - then preindex up by immediate value)
                        {
                            inst.gip_ins_subclass = gip_ins_subclass_memory_byte | gip_ins_subclass_memory_up | gip_ins_subclass_memory_preindex;
                            inst.immediate[4;0] = 0;
                            inst.rm_is_imm = 1;
                            inst.gip_ins_rm.type = gip_ins_r_type_none;
                        }
                        case gip_native_ins_subclass_memory_word_preindex_up: // Preindex Up Word, immediate of four (unless extended - then preindex up by immediate value)
                        {
                            inst.gip_ins_subclass = gip_ins_subclass_memory_word | gip_ins_subclass_memory_up | gip_ins_subclass_memory_preindex;
                            inst.immediate[4;0] = 4;
                            inst.rm_is_imm = 1;
                            inst.gip_ins_rm.type = gip_ins_r_type_none;
                        }
                        case gip_native_ins_subclass_memory_word_preindex_up_shf: // Preindex Up Word by SHF
                        {
                            inst.gip_ins_subclass = gip_ins_subclass_memory_word | gip_ins_subclass_memory_up | gip_ins_subclass_memory_preindex;
                            inst.gip_ins_rm.type = gip_ins_r_type_internal;
                            inst.gip_ins_rm.r = gip_ins_rnm_int_shf;
                            inst.rm_is_imm = 0;
                        }
                        case gip_native_ins_subclass_memory_word_preindex_down_shf: // Preindex Down Word by SHF
                        {
                            inst.gip_ins_subclass = gip_ins_subclass_memory_word | gip_ins_subclass_memory_down | gip_ins_subclass_memory_preindex;
                            inst.gip_ins_rm.type = gip_ins_r_type_internal;
                            inst.gip_ins_rm.r = gip_ins_rnm_int_shf;
                            inst.rm_is_imm = 0;
                        }
                        case gip_native_ins_subclass_memory_word_postindex_up: // Postindex Up Word, immediate of four (unless extended - then preindex up by immediate value)
                        {
                            inst.gip_ins_subclass = gip_ins_subclass_memory_word | gip_ins_subclass_memory_up | gip_ins_subclass_memory_postindex;
                            inst.immediate[4;0] = 4;
                            inst.rm_is_imm = 1;
                            inst.gip_ins_rm.type = gip_ins_r_type_none;
                        }
                        case gip_native_ins_subclass_memory_word_postindex_down: // Postindex down Word, immediate of four (unless extended - then preindex up by immediate value)
                        {
                            inst.gip_ins_subclass = gip_ins_subclass_memory_word | gip_ins_subclass_memory_down | gip_ins_subclass_memory_postindex;
                            inst.immediate[4;0] = 4;
                            inst.rm_is_imm = 1;
                            inst.gip_ins_rm.type = gip_ins_r_type_none;
                        }
                        }
                        if (extended_immediate!=0)
                        {
                            inst.immediate[28;0] = extended_immediate;
                            inst.immediate[31] = extended_immediate[27];
                            inst.immediate[30] = extended_immediate[27];
                            inst.immediate[29] = extended_immediate[27];
                            inst.immediate[28] = extended_immediate[27];
                        }
                        if (extended_rd.type!=gip_ins_r_type_no_override)
                        {
                            inst.rm_is_imm = 0;
                        }
                    }
                    else // Store - code is STR rm, address_mode(rd)
                    {
                        /*b Decode mode and operation, rm
                         */
                        inst.rm_is_imm = 0;
                        // rm (data to store) defaults to native_mapped_rm
                        // rn (address to store) defaults to native_mapped_rn
                        if (!extended_cmd.extended)
                        {
                            inst.a = 1;
                            inst.s_or_stack = 0;
                            inst.k = 0;
                        }
                        inst.gip_ins_class = gip_ins_class_store;

                        full_switch (ins_subclass_ldst)
                        {
                        case gip_native_ins_subclass_memory_word_noindex: // Postindex Up Word, no setting accumulator ; should not extend with rd set to something!
                        {
                            inst.a = 0;
                            inst.gip_ins_subclass = gip_ins_subclass_memory_word | gip_ins_subclass_memory_up | gip_ins_subclass_memory_postindex;
                            inst.gip_ins_rd.type = gip_ins_r_type_none; // No writeback
                        }
                        case gip_native_ins_subclass_memory_half_noindex: // Postindex Up Half, no setting accumulator ; should not extend with rd set to something!
                        {
                            inst.a = 0;
                            inst.gip_ins_subclass = gip_ins_subclass_memory_half | gip_ins_subclass_memory_up | gip_ins_subclass_memory_postindex;
                            inst.gip_ins_rd.type = gip_ins_r_type_none; // No writeback
                        }
                        case gip_native_ins_subclass_memory_byte_noindex: // Postindex Up Byte, no setting accumulator ; should not extend with rd set to something!
                        {
                            inst.a = 0;
                            inst.gip_ins_subclass = gip_ins_subclass_memory_byte | gip_ins_subclass_memory_up | gip_ins_subclass_memory_postindex;
                            inst.gip_ins_rd.type = gip_ins_r_type_none; // No writeback
                        }
                        case gip_native_ins_subclass_memory_word_preindex_up: // Preindex Up Word with writeback
                        {
                            inst.gip_ins_subclass = gip_ins_subclass_memory_word | gip_ins_subclass_memory_up | gip_ins_subclass_memory_preindex;
                            if (extended_rd.type==gip_ins_r_type_no_override)
                            {
                                inst.gip_ins_rd = inst.gip_ins_rn;
                            }
                        }
                        case gip_native_ins_subclass_memory_word_preindex_up_shf: // Preindex Up Word by SHF
                        {
                            inst.gip_ins_subclass = gip_ins_subclass_memory_word | gip_ins_subclass_memory_up | gip_ins_subclass_memory_preindex;
                            inst.p_or_offset_is_shift = 1;
                            inst.gip_ins_rd.type = gip_ins_r_type_none; // No writeback
                        }
                        case gip_native_ins_subclass_memory_word_preindex_down_shf: // Preindex Down Word by SHF
                        {
                            inst.gip_ins_subclass = gip_ins_subclass_memory_word | gip_ins_subclass_memory_down | gip_ins_subclass_memory_preindex;
                            inst.p_or_offset_is_shift = 1;
                            inst.gip_ins_rd.type = gip_ins_r_type_none; // No writeback
                        }
                        case gip_native_ins_subclass_memory_word_postindex_up: // Postindex Up Word
                        {
                            inst.gip_ins_subclass = gip_ins_subclass_memory_word | gip_ins_subclass_memory_up | gip_ins_subclass_memory_postindex;
                            if (extended_rd.type==gip_ins_r_type_no_override)
                            {
                                inst.gip_ins_rd = inst.gip_ins_rn;
                            }
                        }
                        case gip_native_ins_subclass_memory_word_postindex_down: // Postindex down Word
                        {
                            inst.gip_ins_subclass = gip_ins_subclass_memory_word | gip_ins_subclass_memory_down | gip_ins_subclass_memory_postindex;
                            if (extended_rd.type==gip_ins_r_type_no_override)
                            {
                                inst.gip_ins_rd = inst.gip_ins_rn;
                            }
                        }
                        }
                    }
                    /*b Tidy up - common stuff for ldr and str
                     */
                    if (extended_cmd.extended)
                    {
                        if (extended_cmd.op[0])
                        {
                            inst.k = special_repeat_count[4;0];
                        }
                        else
                        {
                            inst.k = extended_cmd.burst;
                        }
                        if (extended_cmd.op[1])
                        {
                            inst.gip_ins_subclass = inst.gip_ins_subclass &~ gip_ins_subclass_memory_index;
                            inst.gip_ins_subclass = inst.gip_ins_subclass | gip_ins_subclass_memory_postindex;
                        }
                        else
                        {
                            inst.gip_ins_subclass = inst.gip_ins_subclass &~ gip_ins_subclass_memory_index;
                            inst.gip_ins_subclass = inst.gip_ins_subclass | gip_ins_subclass_memory_preindex;
                        }
                    }
                    next_extended_cmd.burst = (inst.k==0)?0:(inst.k-1);
                    inst.f = native_mapped_rd_is_pc;
                    inst.valid = 1;
                }
                /*b Special instructions
                 */
                case gip_native_ins_class_special:
                {
                    if (!opcode[0]) // RestartAt instruction
                    {
                        inst.gip_ins_class = gip_ins_class_arith;
                        inst.gip_ins_subclass = gip_ins_subclass_arith_add;
                        inst.a = 0;
                        inst.s_or_stack = 0;
                        inst.p_or_offset_is_shift = 0;
                        inst.f = 0;
                        inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc};
                        inst.gip_ins_rd = {type=gip_ins_r_type_special, r=gip_special_reg_thread_pc};
                        inst.rm_is_imm = 1;
                        inst.immediate = native_mapped_branch_offset;

                        inst.valid = 1;
                        pc_op = gip_pc_op_sequential;
                    }
                    else // block, restart semaphores, restart mode
                    {
                        full_switch (opcode[3;9])
                            {
                            case 0: // restart data
                            {
                                inst.gip_ins_class = gip_ins_class_logic;
                                inst.gip_ins_subclass = gip_ins_subclass_logic_mov;
                                inst.a = 0;
                                inst.s_or_stack = 0;
                                inst.p_or_offset_is_shift = 0;
                                inst.f = 0;
                                inst.gip_ins_rd = {type=gip_ins_r_type_special, r=gip_special_reg_thread_data};
                                inst.rm_is_imm = 1;
                                inst.immediate[8;0] = opcode[8;1];

                                inst.valid = 1;
                                pc_op = gip_pc_op_sequential;
                            }
                            case 1: // block/atomic/deschedule
                            {
                                inst.gip_ins_class = gip_ins_class_logic;
                                inst.gip_ins_subclass = gip_ins_subclass_logic_mov;
                                inst.a = 0;
                                inst.s_or_stack = 0;
                                inst.p_or_offset_is_shift = 0;
                                inst.f = 0;
                                if (opcode[7])
                                {
                                    inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_rnm_int_block_all};
                                }
                                else
                                {
                                    inst.gip_ins_rn.type=gip_ins_r_type_none;
                                }
                                inst.gip_ins_rm.type=gip_ins_r_type_none;
                                inst.gip_ins_rd.type=gip_ins_r_type_none;
                                if (opcode[8])
                                {
                                    inst.tag = 1;
                                    inst.f = 1;
                                }
                                inst.valid = 1;
                                pc_op = gip_pc_op_sequential;
                                next_atomic = opcode[6;1];
                            }
                            case 2:
                            {
                                inst.valid = 0;
                            }
                            case 3:
                            {
                                inst.valid = 0;
                            }
                            case 4:
                            {
                                inst.valid = 0;
                            }
                            case 5:
                            {
                                inst.valid = 0;
                            }
                            case 6:
                            {
                                inst.valid = 0;
                            }
                            case 7:
                            {
                                inst.valid = 0;
                            }
                            }
                    }
                }
                /*b Branch instructions
                 */
                case gip_native_ins_class_branch:
                {
                    /*b Unconditional - build an unconditional reset of condition passed - i.e. AND pc, #0 -> EQ
                     */
                    if (!in_conditional_shadow)
                    {
                        inst.gip_ins_class = gip_ins_class_logic;
                        inst.gip_ins_subclass = gip_ins_subclass_logic_and;
                        inst.a = 0;
                        inst.s_or_stack = 0;
                        inst.p_or_offset_is_shift = 0;
                        inst.f = 0;
                        inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc};
                        inst.gip_ins_rd = {type=gip_ins_r_type_internal, r=gip_ins_rd_int_eq};
                        inst.rm_is_imm = 1;
                        inst.gip_ins_rm.type = gip_ins_r_type_none;
                        inst.immediate = 0;
                        if (branch_delay_slot)
                        {
                            //next_delay_pc =pc+8+native_mapped_branch_offset; always is
                            pc_op = gip_pc_op_delayed_branch; // pc+8+native_mapped_branch_offset;
                            //next_follow_delay_pc = 1;
                            //next_in_delay_slot = 1;
                        }
                        else
                        {
                            pc_op = gip_pc_op_branch; // pc+8+native_mapped_branch_offset;
                        }
                    }
                    /*b Build a conditional flushing instruction (ADD<cc>F pc, #offset), mark next instruction as delayed if required
                     */
                    else
                    {
                        inst.gip_ins_class = gip_ins_class_arith;
                        inst.gip_ins_subclass = gip_ins_subclass_arith_add;
                        inst.a = 0;
                        inst.s_or_stack = 0;
                        inst.p_or_offset_is_shift = 0;
                        inst.f = 1;
                        inst.gip_ins_rn = {type=gip_ins_r_type_internal, r=gip_ins_r_int_pc};
                        inst.gip_ins_rd = {type=gip_ins_r_type_internal, r=gip_ins_rd_int_eq};
                        inst.rm_is_imm = 1;
                        inst.gip_ins_rm.type = gip_ins_r_type_none;
                        inst.immediate = native_mapped_branch_offset;
                        //next_in_delay_slot = branch_delay_slot;
                    }
                    inst.valid = 1;
                }
                /*b Done all instructions
                 */
                default:
                {
                    pc_op = gip_pc_op_sequential;
                }
                }
        }

    /*b Done
     */
}
