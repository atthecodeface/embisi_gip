/*a Includes
 */
include "gip.h"
include "gip_internal.h"

/*a Modules
 */
module gip_alu_logical_op( input t_gip_word op_a,
                           input t_gip_word op_b,
                           input t_gip_logic_op logic_op,
                           input bit z_in,
                           input bit n_in,
                           input bit c_in,
                           input bit v_in,
                           output t_gip_word result,
                           output bit z,
                           output bit n )
"
This module implements the logical operations for the GIP
"
{
    comb t_gip_word anded;
    comb t_gip_word xored;
    comb bit[8] bit_reversed_byte;
    comb t_gip_word byte_reversed;
    comb bit[6] counted;
    comb bit[6] counted_a;
    comb bit[8] anded_a;
    comb bit[6] counted_b;
    comb bit[8] anded_b;
    comb bit[6] counted_c;
    comb bit[8] anded_c;
    comb bit[6] counted_d;
    comb bit[8] anded_d;
    comb bit[8] first_bit_byte;
    comb bit[5] first_bit_number;
   
    /*b First steps
     */
    first_steps "First steps of operation":
        {
            anded = op_a & op_b;
            xored = op_a ^ op_b;

            for (i; 8)
            {
                bit_reversed_byte[7-i] = op_b[i];
            }

            byte_reversed[8;24] = op_b[8; 0];
            byte_reversed[8;16] = op_b[8; 8];
            byte_reversed[8; 8] = op_b[8;16];
            byte_reversed[8; 0] = op_b[8;24];
        }

    /*b Count bits
     */
    count_bits "Count bits in anded[]":
        {
            counted_a = 0;
            anded_a = anded[8;0];
            for (i; 8)
            {
                if (anded_a[i])
                {
                    counted_a = counted_a + 1;
                }
            }

            counted_b = 0;
            anded_b = anded[8;8];
            for (i; 8)
            {
                if (anded_b[i])
                {
                    counted_b = counted_b + 1;
                }
            }

            counted_c = 0;
            anded_c = anded[8;16];
            for (i; 8)
            {
                if (anded_c[i])
                {
                    counted_c = counted_c + 1;
                }
            }

            counted_d = 0;
            anded_d = anded[8;24];
            for (i; 8)
            {
                if (anded_d[i])
                {
                    counted_d = counted_d + 1;
                }
            }
            counted = counted_a + counted_b + counted_c + counted_d;

        }

    /*b Find first bit set
     */
    first_bit "Determine first bit set (from top) in xored - zero for none as well as bit 0":
        {
            first_bit_number = 0;
            if (xored[8;24]!=0)
            {
                first_bit_byte = xored[8;24];
                first_bit_number[2;3] = 3;
            }
            elsif (xored[8;16]!=0)
            {
                first_bit_byte = xored[8;16];
                first_bit_number[2;3] = 2;
            }
            elsif (xored[8;8]!=0)
            {
                first_bit_byte = xored[8;8];
                first_bit_number[2;3] = 1;
            }
            else
            {
                first_bit_byte = xored[8;0];
                first_bit_number[2;3] = 0;
            }
            if (first_bit_byte[4;4] != 0)
            {
                if (first_bit_byte[7]) { first_bit_number[3;0] = 7; }
                elsif (first_bit_byte[6]) { first_bit_number[3;0] = 6; }
                elsif (first_bit_byte[5]) { first_bit_number[3;0] = 5; }
                else { first_bit_number[3;0] = 4; }
            }
            else
            {
                if (first_bit_byte[3]) { first_bit_number[3;0] = 3; }
                elsif (first_bit_byte[2]) { first_bit_number[3;0] = 2; }
                elsif (first_bit_byte[1]) { first_bit_number[3;0] = 1; }
                else { first_bit_number[3;0] = 0; }
            }
        }

    /*b Final result
     */
    final_result "Final result selection/operation":
        {
            result = 0;
            part_switch (logic_op)
                {
                case gip_logic_op_mov: { result =          op_b; }
                case gip_logic_op_mvn: { result =         ~op_b; }
                case gip_logic_op_and: { result =  op_a &  op_b; }
                case gip_logic_op_or:  { result =  op_a |  op_b; }
                case gip_logic_op_xor: { result =  op_a ^  op_b; }
                case gip_logic_op_bic: { result =  op_a & ~op_b; }
                case gip_logic_op_orn: { result =  op_a | ~op_b; }
                case gip_logic_op_and_xor: { result =  anded ^  op_b; }
                case gip_logic_op_and_cnt: { result[6;0] = counted; }
                case gip_logic_op_xor_first: { result[5;0] = first_bit_number; }
                case gip_logic_op_bit_reverse: { result = op_b; result[8;0] = bit_reversed_byte; }
                case gip_logic_op_byte_reverse: { result = byte_reversed; }
                case gip_logic_op_read_flags: { result[0] = z_in; result[1] = n_in; result[2] = c_in; result[3] = v_in; }
                }
            z = (result==0);
            n = result[31];
        }

    /*b Done
     */
}
