/*a Includes
 */
include "postbus.h"

/*a Types
 */
/*t t_arb_fsm
 */
typedef fsm
{
    arb_fsm_idle;
    arb_fsm_src_0;
    arb_fsm_src_1;
    arb_fsm_src_2;
    arb_fsm_src_3;
} t_arb_fsm;

/*t t_buf_fsm
 */
typedef fsm
{
    buf_fsm_idle; // Buffers both empty - fill 0 first
    buf_fsm_0_rdy; // Buffer 0 is full, present it to target
    buf_fsm_0_rdy_1_pend; // Buffer 0 is full, 1 also (to follow 0); present 0 to target
    buf_fsm_1_rdy; // Buffer 1 is full, present it to target
    buf_fsm_1_rdy_0_pend; // Buffer 1 is full, 0 also (to follow 1); present 1 to target
    buf_fsm_wait; // No buffers full, but in middle of transaction
} t_buf_fsm;

typedef struct
{
    t_postbus_data data;
    bit first;
    bit last;
} t_buf_data;
/*a postbus_register_demux module
 */
module postbus_register_demux( clock int_clock, input bit int_reset,
                               input t_postbus_type src_type, input t_postbus_data src_data, output t_postbus_ack src_ack,
                               input t_postbus_ack tgt_ack_0, output t_postbus_type tgt_type_0,
                               input t_postbus_ack tgt_ack_1, output t_postbus_type tgt_type_1,
                               input t_postbus_ack tgt_ack_2, output t_postbus_type tgt_type_2,
                               input t_postbus_ack tgt_ack_3, output t_postbus_type tgt_type_3,
                               output t_postbus_data tgt_data 
    )
    "This is a 1-to-4 dual-word buffer register postbus demultiplexer.
    It should be driven by an n-to-1 multiplexer.
    It should drive a number of final combinatorial p-to-q postbus multiplexers."
{
    /*b State and combinatorials
     */
    default clock rising int_clock;
    default reset active_high int_reset;

    clocked t_buf_fsm buf_state = buf_fsm_idle;
    comb t_buf_fsm next_buf_state "Next state of buffer FSM";

    clocked t_buf_data[2] buffer = { { data=0,first=0,last=0 }, { data=0,first=0,last=0 }};

    clocked bit[2] last_target = 0;
    comb bit[2] selected_target;

    comb bit src_first;
    comb bit src_last;

    comb bit[2] buffer_write_enable;
    comb bit buffer_read;

    comb t_postbus_type tgt_type;
    comb t_postbus_ack tgt_ack;

    /*b Buffer state FSM - src_first, src_last
     */
    src_first_last "Determine first/last indications for the current source presented word":
        {
            src_first = 0;
            src_last = 0;
            part_switch (src_type)
            {
            case postbus_word_type_start:
            {
                src_first = 1;
                src_last = src_data[0];
            }
            case postbus_word_type_last:
            {
                src_last = 1;
            }
            }
        }

    /*b Buffer buf_state FSM - buf_state, next_buf_state, buffer_write_enable, src_ack, buffer_read
     */
    buffer_fsm "Buffer state FSM - move on if data is given or taken away":
        {
            next_buf_state = buf_state;
            buffer_write_enable = 0;
            src_ack = 0;
            buffer_read = 0;
            full_switch (buf_state)
                {
                case buf_fsm_idle:
                {
                    src_ack = 1;
                    if (src_type==postbus_word_type_start)
                    {
                        next_buf_state = buf_fsm_0_rdy;
                        buffer_write_enable[0] = 1;
                    };
                }
                case buf_fsm_0_rdy:
                {
                    src_ack = 1;
                    if (src_type!=postbus_word_type_idle)
                    {
                        if (tgt_ack)
                        {
                            next_buf_state = buf_fsm_1_rdy;
                        }
                        else
                        {
                            next_buf_state = buf_fsm_0_rdy_1_pend;
                        }
                        buffer_write_enable[1] = 1;
                    }
                }
                case buf_fsm_1_rdy:
                {
                    src_ack = 1;
                    buffer_read = 1;
                    if (src_type!=postbus_word_type_idle)
                    {
                        if (tgt_ack)
                        {
                            next_buf_state = buf_fsm_0_rdy;
                        }
                        else
                        {
                            next_buf_state = buf_fsm_1_rdy_0_pend;
                        }
                        buffer_write_enable[0] = 1;
                    }
                }
                case buf_fsm_0_rdy_1_pend:
                {
                    if (tgt_ack)
                    {
                        next_buf_state = buf_fsm_1_rdy;
                    }
                }
                case buf_fsm_1_rdy_0_pend:
                {
                    buffer_read = 1;
                    if (tgt_ack)
                    {
                        next_buf_state = buf_fsm_0_rdy;
                    }
                }
                }
            buf_state <= next_buf_state;
        }

    /*b Output select for target type, target data - tgt_type, tgt_data
     */
    target_type_output "Output select for target type":
        {
            tgt_type = postbus_word_type_data;
            if (buffer[buffer_read].last)
            {
                tgt_type = postbus_word_type_start;
            }
            if (buffer[buffer_read].first)
            {
                tgt_type = postbus_word_type_last;
            }
            if (buf_state==buf_fsm_idle)
            {
                tgt_type = postbus_word_type_idle;
            }
            tgt_data = buffer[buffer_read].data;
        }

    /*b Multiplexer/Demultiplexer for selected target - tgt_type_*, tgt_ack
     */
    target_mux_demux "Multiplexer/Demultiplexer for selected target":
        {
            tgt_type_0 = postbus_word_type_idle;
            tgt_type_1 = postbus_word_type_idle;
            tgt_type_2 = postbus_word_type_idle;
            tgt_type_3 = postbus_word_type_idle;
            full_switch (selected_target)
            {
            case 0: {tgt_type_0 = tgt_type; tgt_ack=tgt_ack_0;}
            case 1: {tgt_type_1 = tgt_type; tgt_ack=tgt_ack_1;}
            case 2: {tgt_type_2 = tgt_type; tgt_ack=tgt_ack_2;}
            case 3: {tgt_type_3 = tgt_type; tgt_ack=tgt_ack_3;}
            }
        }

    /*b Selected target - selected_target, last_target
     */
    selected_target "Selected target and last_target register":
        {
            // selected_target comes out of current read buffer if that has a first word; else out of last_target_register
            // last_target_register is stored every time the current read buffer has a first word
            selected_target = last_target;
            if (buffer[buffer_read].first)
            {
                selected_target = buffer[buffer_read].data[2;1];
                last_target <= selected_target;
            }
        }

    /*b Data buffer - buffer
     */
    data_buffer "Data buffer":
        {
            for ( i; 2 )
            {
                if (buffer_write_enable[i])
                {
                    if (i==0)
                    {
                        buffer[0].data <= src_data;
                    }
                    else
                    {
                        buffer[1].data <= src_data;
                    }
                    buffer[i].first <= src_first;
                    buffer[i].last <= src_last;
                }
            }
        }

    /*b Done
     */
}
