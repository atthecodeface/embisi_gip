/*a Includes
 */
include "gip.h"
include "gip_internal.h"

/*a Modules
 */
module gip_alu_logical_op( input t_gip_word op_a,
                           input t_gip_word op_b,
                           input t_gip_logic_op logic_op,
                           input bit z_in,
                           input bit n_in,
                           input bit c_in,
                           input bit v_in,
                           output t_gip_word result,
                           output bit z,
                           output bit n )
"
This module implements the logical operations for the GIP
"
{
    //comb t_gip_word anded;
    //comb t_gip_word xored;
    //comb bit[8] bit_reversed_byte;
    //comb t_gip_word byte_reversed;
    //comb bit[6] counted;
    //comb bit[6] counted_a;
    //comb bit[8] anded_a;
    //comb bit[6] counted_b;
    //comb bit[8] anded_b;
    //comb bit[6] counted_c;
    //comb bit[8] anded_c;
    //comb bit[6] counted_d;
    //comb bit[8] anded_d;
    //comb bit[8] first_bit_byte;
    //comb bit[5] first_bit_number;
   
    /*b Final result
     */
    final_result "Final result selection/operation":
        {
            result = 0;
            part_switch (logic_op)
                {
                case gip_logic_op_mov: { result =          op_b; }
                case gip_logic_op_mvn: { result =         ~op_b; }
                case gip_logic_op_and: { result =  op_a &  op_b; }
                case gip_logic_op_or:  { result =  op_a |  op_b; }
                case gip_logic_op_xor: { result =  op_a ^  op_b; }
                case gip_logic_op_bic: { result =  op_a & ~op_b; }
                case gip_logic_op_orn: { result =  op_a | ~op_b; }
                    //case gip_logic_op_and_xor: { result =  anded ^  op_b; }
                    //case gip_logic_op_and_cnt: { result[6;0] = counted; }
                    //case gip_logic_op_xor_first: { result[5;0] = first_bit_number; }
                    //case gip_logic_op_bit_reverse: { result = op_b; result[8;0] = bit_reversed_byte; }
                    //case gip_logic_op_byte_reverse: { result = byte_reversed; }
                case gip_logic_op_read_flags: { result[0] = z_in; result[1] = n_in; result[2] = c_in; result[3] = v_in; }
                }
            z = (result==0);
            n = result[31];
        }

    /*b Done
     */
}
