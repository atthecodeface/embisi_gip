/*a To do
  Block on memory busy, memory transaction in progress
  Block on rfw busy, rfw required
 */

/*a Includes
 */
include "gip.h"
include "gip_internal.h"
include "gip_alu.h"

/*a Types
 */
/*t t_gip_alu_flags
 */
typedef struct
{
    bit z;
    bit n;
    bit c;
    bit v;
    bit p;
    bit cp;
    bit old_cp;
} t_gip_alu_flags;

/*a Module
 */
module gip_alu( clock gip_clock,
                input bit gip_reset,

                input t_gip_instruction_rf rfr_inst,
                input t_gip_word rf_read_port_0,
                input t_gip_word rf_read_port_1,

                output t_gip_instruction_rf alu_inst,

                input bit rfw_accepting_alu_rd,
                input bit mem_alu_busy,
                input bit alu_accepting_rfr_instruction,
                output bit alu_accepting_rfr_instruction_always,
                output bit alu_accepting_rfr_instruction_if_mem_does,
                output bit alu_accepting_rfr_instruction_if_rfw_does,

                output t_gip_ins_r alu_rd,
                output bit alu_use_shifter,
                output t_gip_word alu_arith_logic_result,
                output t_gip_word alu_shifter_result,

                output t_gip_mem_op alu_mem_op,
                output t_gip_mem_options alu_mem_options,
                output t_gip_ins_r alu_mem_rd,
                output t_gip_word alu_mem_address,
                output t_gip_word alu_mem_write_data,
                output bit[4] alu_mem_burst,

                input bit special_cp_trail_2,

                output bit gip_pipeline_flush,
                output bit[2] gip_pipeline_tag,
                output bit gip_pipeline_executing
    )
{
    /*b Default clock and reset
     */
    default clock gip_clock;
    default reset gip_reset;

    comb bit writes_conditional;
    comb bit conditional_result;

    comb t_gip_word alu_op1;
    comb t_gip_word alu_op2;

    comb bit set_zcvn;
    comb bit set_p;
    comb bit set_acc;
    comb t_gip_arith_op gip_arith_op;
    comb t_gip_logic_op gip_logic_op;
    comb t_gip_shift_op gip_shift_op;
    comb t_gip_word alu_constant;

    comb bit shf_carry_in;
    comb t_gip_word shf_value_in;
    comb bit[8] shf_amount_in;

    net bit shf_carry;
    net t_gip_word shf_result;

    net bit arith_z;
    net bit arith_n;
    net bit arith_c;
    net bit arith_v;
    net t_gip_word arith_result;
    net bit shf_carry_override_value;
    net bit shf_carry_override;
    comb bit shf_carry_overridden;

    net bit logic_z;
    net bit logic_n;
    net t_gip_word logic_result;

    comb bit condition_passed;

    clocked t_gip_instruction_rf alu_inst =
        {
            valid=0,
            gip_ins_class=gip_ins_class_logic,
            gip_ins_subclass=gip_ins_subclass_logic_mov,
            gip_ins_cc=gip_ins_cc_always,
            gip_ins_rd={type=gip_ins_r_type_register,r=0},
            gip_ins_rn={type=gip_ins_r_type_register,r=0},
            gip_ins_rm={type=gip_ins_r_type_register,r=0},
            rm_is_imm = 0,
            immediate=0,
            k=0,
            a=0,
            f=0,
            s_or_stack=0,
            p_or_offset_is_shift=0,
            d=0,
            pc=0,
            tag=0
        };
    clocked bit first_cycle_of_instruction = 0;

    clocked t_gip_word alu_a_in=0;
    clocked t_gip_word alu_b_in=0;
    clocked t_gip_word shf=0;
    clocked t_gip_word acc=0;
    clocked t_gip_alu_flags flags = {z=0, n=0, v=0, c=0, p=0, cp=0, old_cp=0};

    comb t_gip_alu_flags next_flags;
    comb t_gip_word next_shf;
    comb t_gip_word next_acc;

    comb t_gip_alu_op1_src alu_op1_src;
    comb t_gip_alu_op2_src alu_op2_src;

    /*b Evaluate condition associated with the instruction - simultaneous with ALU stage, blocks all results from instruction if it fails; depends directly on state
     */
    condition_passed "Evaluate condition associated with the instruction - simultaneous with ALU stage, blocks all results from instruction if it fails":
        {
            condition_passed = 0;
            if (alu_inst.valid)
            {
                part_switch (alu_inst.gip_ins_cc )
                    {
                    case gip_ins_cc_eq: { condition_passed = flags.z; }
                    case gip_ins_cc_ne: { condition_passed = !flags.z; }
                    case gip_ins_cc_cs: { condition_passed = flags.c; }
                    case gip_ins_cc_cc: { condition_passed = !flags.c; }
                    case gip_ins_cc_mi: { condition_passed = flags.n; }
                    case gip_ins_cc_pl: { condition_passed = !flags.n; }
                    case gip_ins_cc_vs: { condition_passed = flags.v; }
                    case gip_ins_cc_vc: { condition_passed = !flags.v; }
                    case gip_ins_cc_hi: { condition_passed = flags.c && !flags.z; }
                    case gip_ins_cc_ls: { condition_passed = !flags.c || flags.z; }
                    case gip_ins_cc_ge: { condition_passed = (!flags.n && !flags.v) || (flags.n && flags.v); }
                    case gip_ins_cc_lt: { condition_passed = (!flags.n && flags.v) || (flags.n && !flags.v); }
                    case gip_ins_cc_gt: { condition_passed = ((!flags.n && !flags.v) || (flags.n && flags.v)) && !flags.z; }
                    case gip_ins_cc_le: { condition_passed = ((!flags.n && flags.v) || (flags.n && !flags.v)) || flags.z; }
                    case gip_ins_cc_always: { condition_passed = 1; }
                    case gip_ins_cc_cp: { condition_passed = special_cp_trail_2 ? (flags.cp && flags.old_cp) : flags.cp; }
                    }
            }
        }

    /*b Determine which flags and accumulator to set, and the ALU operation; depends on state (except shf_value and shf_value, which depends on alu_op1/2)
     */
    determine_operation "Determine operation":
        {
            alu_use_shifter = 0;
            gip_arith_op = gip_arith_op_add;
            gip_logic_op = gip_logic_op_mov;
            gip_shift_op = gip_shift_op_lsl;
            shf_carry_in = 0;
            shf_value_in = alu_op1;
            shf_amount_in = 0;
            part_switch (alu_inst.gip_ins_class)
            {
            case gip_ins_class_arith:
            {
                part_switch (alu_inst.gip_ins_subclass)
                    {
                    case gip_ins_subclass_arith_add:  {gip_arith_op = gip_arith_op_add;}
                    case gip_ins_subclass_arith_adc:  {gip_arith_op = gip_arith_op_adc;}
                    case gip_ins_subclass_arith_sub:  {gip_arith_op = gip_arith_op_sub;}
                    case gip_ins_subclass_arith_sbc:  {gip_arith_op = gip_arith_op_sbc;}
                    case gip_ins_subclass_arith_rsb:  {gip_arith_op = gip_arith_op_rsub;}
                    case gip_ins_subclass_arith_rsc:  {gip_arith_op = gip_arith_op_rsbc;}
                    case gip_ins_subclass_arith_init:
                    {
                        gip_arith_op = gip_arith_op_init;
                        shf_carry_in = 0;
                        gip_shift_op = gip_shift_op_lsr;
                        shf_value_in = alu_op1;
                        shf_amount_in = 0;
                    }
                    case gip_ins_subclass_arith_mla:
                    {
                        gip_arith_op = gip_arith_op_mla;
                        shf_carry_in = flags.c;
                        gip_shift_op = gip_shift_op_lsr;
                        shf_value_in = shf;
                        shf_amount_in = 2;
                    }
                    case gip_ins_subclass_arith_mlb:
                    {
                        gip_arith_op = gip_arith_op_mlb;
                        shf_carry_in = flags.c;
                        gip_shift_op = gip_shift_op_lsr;
                        shf_value_in = shf;
                        shf_amount_in = 2;
                    }
                    case gip_ins_subclass_arith_write_flags:  {gip_arith_op = gip_arith_op_write_flags;}
                    }
            }
            case gip_ins_class_logic:
            {
                part_switch (alu_inst.gip_ins_subclass)
                    {
                    case gip_ins_subclass_logic_and:  {gip_logic_op = gip_logic_op_and;}
                    case gip_ins_subclass_logic_or:   {gip_logic_op = gip_logic_op_or;}
                    case gip_ins_subclass_logic_xor:  {gip_logic_op = gip_logic_op_xor;}
                    case gip_ins_subclass_logic_bic:  {gip_logic_op = gip_logic_op_bic;}
                    case gip_ins_subclass_logic_orn:  {gip_logic_op = gip_logic_op_orn;}
                    case gip_ins_subclass_logic_mov:  {gip_logic_op = gip_logic_op_mov;}
                    case gip_ins_subclass_logic_mvn:  {gip_logic_op = gip_logic_op_mvn;}
                    case gip_ins_subclass_logic_andcnt:  {gip_logic_op = gip_logic_op_and_cnt;}
                    case gip_ins_subclass_logic_andxor:  {gip_logic_op = gip_logic_op_and_xor;}
                    case gip_ins_subclass_logic_xorfirst:  {gip_logic_op = gip_logic_op_xor_first;}
                    case gip_ins_subclass_logic_bitreverse:  {gip_logic_op = gip_logic_op_bit_reverse;}
                    case gip_ins_subclass_logic_bytereverse:  {gip_logic_op = gip_logic_op_byte_reverse;}
                    case gip_ins_subclass_logic_read_flags:  {gip_logic_op = gip_logic_op_read_flags;}
                    }
            }
            case gip_ins_class_shift:
            {
                alu_use_shifter = 1;
                part_switch (alu_inst.gip_ins_subclass)
                    {
                    case gip_ins_subclass_shift_lsl:
                    {
                        shf_carry_in = flags.c;
                        gip_shift_op = gip_shift_op_lsl;
                        shf_value_in = alu_op1;
                        shf_amount_in = alu_op2[8;0];
                    }
                    case gip_ins_subclass_shift_lsr:
                    {
                        shf_carry_in = flags.c;
                        gip_shift_op = gip_shift_op_lsr;
                        shf_value_in = alu_op1;
                        shf_amount_in = alu_op2[8;0];
                    }
                    case gip_ins_subclass_shift_asr:
                    {
                        shf_carry_in = flags.c;
                        gip_shift_op = gip_shift_op_asr;
                        shf_value_in = alu_op1;
                        shf_amount_in = alu_op2[8;0];
                    }
                    case gip_ins_subclass_shift_ror:
                    {
                        shf_carry_in = flags.c;
                        gip_shift_op = gip_shift_op_ror;
                        shf_value_in = alu_op1;
                        shf_amount_in = alu_op2[8;0];
                    }
                    case gip_ins_subclass_shift_ror33:
                    {
                        shf_carry_in = flags.c;
                        gip_shift_op = gip_shift_op_rrx;
                        shf_value_in = alu_op1;
                        shf_amount_in = alu_op2[8;0];
                    }
                    }
            }
            case gip_ins_class_store:
            case gip_ins_class_load:
            {
                if ((alu_inst.gip_ins_subclass & gip_ins_subclass_memory_dirn)==gip_ins_subclass_memory_up)
                {
                    gip_arith_op = gip_arith_op_add;
                }
                else
                {
                    gip_arith_op = gip_arith_op_sub;
                }
            }
            }
        }

    /*b Determine inputs to the shifter and ALU; depends on state, but 32-bit muxes required to get alu_op1/2
     */
    input_determination "Determine inputs to the shifter and ALU":
    {
        alu_op1_src = gip_alu_op1_src_a_in;
        if ( (alu_inst.gip_ins_rn.type == gip_ins_r_type_internal) &&
             (alu_inst.gip_ins_rn.r    == gip_ins_rnm_int_acc) )
        {
            alu_op1_src = gip_alu_op1_src_acc;
        }

        alu_op2_src = gip_alu_op2_src_b_in;
        alu_constant = 0;
        if (!alu_inst.rm_is_imm)
        {
            if ( (alu_inst.gip_ins_rm.type == gip_ins_r_type_internal) &&
                 (alu_inst.gip_ins_rm.r    == gip_ins_rnm_int_acc) )
            {
                alu_op2_src = gip_alu_op2_src_acc;
            }
            if ( (alu_inst.gip_ins_rm.type == gip_ins_r_type_internal) &&
                 (alu_inst.gip_ins_rm.r    == gip_ins_rnm_int_shf) )
            {
                alu_op2_src = gip_alu_op2_src_shf;
            }

            if (alu_inst.gip_ins_class == gip_ins_class_store )
            {
                part_switch (alu_inst.gip_ins_subclass[2;0])
                {
                case gip_ins_subclass_memory_word: { alu_constant = 4; }
                case gip_ins_subclass_memory_half: { alu_constant = 2; }
                case gip_ins_subclass_memory_byte: { alu_constant = 1; }
                }
                if (alu_inst.p_or_offset_is_shift)
                {
                    alu_op2_src = gip_alu_op2_src_shf;
                }
                else
                {
                    alu_op2_src = gip_alu_op2_src_constant;
                }
            }
        }

        alu_op1 = acc;
        alu_op2 = acc;
        part_switch (alu_op1_src)
            {
            case gip_alu_op1_src_a_in: { alu_op1 = alu_a_in; }
            case gip_alu_op1_src_acc:  { alu_op1 = acc; }
            }
        full_switch (alu_op2_src)
            {
            case gip_alu_op2_src_b_in: { alu_op2 = alu_b_in; }
            case gip_alu_op2_src_acc:  { alu_op2 = acc; }
            case gip_alu_op2_src_shf:  { alu_op2 = shf; }
            case gip_alu_op2_src_constant:  { alu_op2 = alu_constant; }
            }
    }

    /*b Perform shifter operation - operates on C, ALU A in, ALU B in: what about accumulator?
     */
    shifter "Perform shifter operation - operates on C, ALU A in, ALU B in: what about accumulator?":
    {
        gip_alu_barrel_shift shift_op( carry_in <= shf_carry_in,
                           gip_shift_op <= gip_shift_op,
                           value <= shf_value_in,
                           amount <= shf_amount_in,
                           result => shf_result,
                           carry_out => shf_carry );
    }

    /*b Perform logical operation - operates on ALU op 1 and ALU op 2
     */
    logical_op "Perform logical operation - operates on ALU op 1 and ALU op 2":
    {
        gip_alu_logical_op logical_op( op_a <= alu_op1,
                                       op_b <= alu_op2,
                                       logic_op <= gip_logic_op,
                                       z_in <= flags.z,
                                       n_in <= flags.n,
                                       c_in <= flags.c,
                                       v_in <= flags.v,
                                       result => logic_result,
                                       z => logic_z,
                                       n => logic_n );
    }

    /*b Perform arithmetic operation - operates on C, ALU op 1 and ALU op 2
     */
    arith_op "Perform arith operation - operates on ALU op 1 and ALU op 2":
    {
        gip_alu_arith_op arith_op( op_a <= alu_op1,
                                   op_b <= alu_op2,
                                   c_in <= flags.c,
                                   p_in <= flags.p,
                                   shf <= shf[2;0],
                                   arith_op <= gip_arith_op,
                                   result => arith_result,
                                   z => arith_z,
                                   n => arith_n,
                                   v => arith_v,
                                   c => arith_c,
                                   shf_carry_override => shf_carry_override,
                                   shf_carry_out => shf_carry_override_value );
    }

    /*b Determine how to set 'cp' and 'old_cp'
     */
    handle_conditional_targets "Determine how to set 'cp' and 'old_cp' with conditional targets":
        {
            writes_conditional = 0;
            conditional_result = 0;
            if (alu_inst.gip_ins_rd.type == gip_ins_r_type_internal) 
            {
                part_switch (alu_inst.gip_ins_rd.r)
                    {
                    case gip_ins_rd_int_eq:
                    {
                        if (alu_inst.gip_ins_class == gip_ins_class_logic)
                        {
                            conditional_result = logic_z;
                        }
                        else
                        {
                            conditional_result = arith_z;
                        }
                        writes_conditional = 1;
                    }
                    case gip_ins_rd_int_ne:
                    {
                        if (alu_inst.gip_ins_class == gip_ins_class_logic)
                        {
                            conditional_result = !logic_z;
                        }
                        else
                        {
                            conditional_result = !arith_z;
                        }
                        writes_conditional = 1;
                    }
                    case gip_ins_rd_int_cs:
                    {
                        conditional_result = arith_c;
                        writes_conditional = 1;
                    }
                    case gip_ins_rd_int_cc:
                    {
                        conditional_result = !arith_c;
                        writes_conditional = 1;
                    }
                    case gip_ins_rd_int_hi:
                    {
                        conditional_result = arith_c && !arith_z;
                        writes_conditional = 1;
                    }
                    case gip_ins_rd_int_ls:
                    {
                        conditional_result = !arith_c || arith_z;
                        writes_conditional = 1;
                    }
                    case gip_ins_rd_int_ge:
                    {
                        conditional_result = (!arith_n && !arith_v) || (arith_n && arith_v);
                        writes_conditional = 1;
                    }
                    case gip_ins_rd_int_lt:
                    {
                        conditional_result = (!arith_n && arith_v) || (arith_n && !arith_v);
                        writes_conditional = 1;
                    }
                    case gip_ins_rd_int_gt:
                    {
                        conditional_result = ((!arith_n && !arith_v) || (arith_n && arith_v)) && !arith_z;
                        writes_conditional = 1;
                    }
                    case gip_ins_rd_int_le:
                    {
                        conditional_result = (!arith_n && arith_v) || (arith_n && !arith_v) || arith_z;
                        writes_conditional = 1;
                    }
                    }
            }
        }

    /*b Determine ALU result, next accumulator, next shifter and next flags
     */
    determine_results "Determine results":
        {
            next_flags = flags;
            next_acc = acc;
            next_shf = shf;
            alu_arith_logic_result = arith_result;
            alu_shifter_result = shf_result;
            set_zcvn = alu_inst.s_or_stack;
            set_p = alu_inst.p_or_offset_is_shift;
            set_acc = alu_inst.a;
            shf_carry_overridden = shf_carry;
            if (shf_carry_override)
            {
                shf_carry_overridden = shf_carry_override_value;
            }
            if (!condition_passed)
            {
                set_acc = 0;
                set_zcvn = 0;
                set_p = 0;
            }
            part_switch (alu_inst.gip_ins_class)
            {
            case gip_ins_class_arith:
            {
                alu_arith_logic_result = arith_result;
                if (set_zcvn)
                {
                    next_flags.z = arith_z;
                    next_flags.c = arith_c;
                    next_flags.v = arith_v;
                    next_flags.n = arith_n;
                }
                if (set_acc)
                {
                    next_acc = arith_result;
                }
                if (set_p)
                {
                    next_shf = shf_result; // Use SHF result if P is not set - this is for init, mla, mlb
                    next_flags.p = shf_carry_overridden; // only for init, mla, mlb
                }
                else
                {
                    next_shf = 0; // Clear SHF if P is set
                }
            }
            case gip_ins_class_logic:
            {
                alu_arith_logic_result = logic_result;
                if (set_p)
                {
                    next_flags.c = flags.p;
                }
                if (set_zcvn)
                {
                    next_flags.z = logic_z;
                    next_flags.n = logic_n;
                }
                if (set_acc)
                {
                    next_acc = logic_result;
                }
            }
            case gip_ins_class_shift:
            {
                if (set_zcvn)
                {
                    next_flags.z = (shf_result==0);
                    next_flags.n = shf_result[31];
                    next_flags.c = shf_carry;
                }
                next_shf = shf_result;
                next_flags.p = shf_carry;
            }
            case gip_ins_class_store:
            case gip_ins_class_load:
            {
                alu_arith_logic_result = arith_result;
                if (set_acc)
                {
                    next_acc = arith_result;
                }
            }
            }
            if (writes_conditional)
            {
                if (condition_passed) // could be first of a sequence, or later on; if first of a sequence, we must set it to our result; if later then condition should be CP for ANDing condition passed
                    // if ANDing (CP is therefore set) and our result is 1, then the next result is 1; if our result is 0, then the next result is zero; so this is the same as the first condition
                {
                    next_flags.cp = conditional_result;
                }
                else // must be later in a sequence; condition ought to have been 'CP', so this means 'state.cp' should be zero already. No reason to make it one.
                {
                    next_flags.cp = 0;
                }
                next_flags.old_cp = 1;
            }
            else
            {
                next_flags.cp = condition_passed;
                next_flags.old_cp = flags.cp;
            }
        }

    /*b Get inputs to memory stage
     */
    memory_stage_inputs "Memory stage inputs":
        {
            if ((alu_inst.gip_ins_subclass & gip_ins_subclass_memory_index)==gip_ins_subclass_memory_preindex)
            {
                alu_mem_address = arith_result;
            }
            else
            {
                alu_mem_address = alu_op1;
            }
            alu_mem_write_data = alu_b_in;
        }

    /*b Determine next Rd for the ALU operation, and memory operation, and if the instruction is blocked - alu_rd, alu_mem_rd, alu_accepting_*
     */
    next_rd_and_blocking "Determine next Rd for the ALU operation, and memory operation, and if the instruction is blocked":
        {
            alu_rd.type = gip_ins_r_type_none;
            alu_rd.r = 0;
            alu_mem_rd.type = gip_ins_r_type_none;
            alu_mem_rd.r = 0;
            alu_mem_op = gip_mem_op_none;
            alu_accepting_rfr_instruction_always = 0;
            alu_accepting_rfr_instruction_if_rfw_does = 0;
            alu_accepting_rfr_instruction_if_mem_does = 0;
            alu_mem_options = gip_mem_options_none;
            if ( alu_inst.s_or_stack ) // indicates stack for memory operations
            {
                alu_mem_options = alu_mem_options | gip_mem_options_stack;
            }
            if (alu_inst.p_or_offset_is_shift ) // indicates signed for memory load operations
            {
                alu_mem_options = alu_mem_options | gip_mem_options_signed; // signed bit should be ignored for stores
            }
            alu_mem_options = alu_mem_options | gip_mem_options_bigendian;
            if (condition_passed) // This is zero if instruction is not valid, so no writeback from invalid instructions!
            {
                part_switch (alu_inst.gip_ins_class)
                {
                case gip_ins_class_arith:
                case gip_ins_class_logic:
                case gip_ins_class_shift:
                {
                    alu_rd = alu_inst.gip_ins_rd;
                    alu_accepting_rfr_instruction_if_rfw_does = 1;
                }
                case gip_ins_class_store:
                {
                    alu_rd = alu_inst.gip_ins_rd;
                    part_switch (alu_inst.gip_ins_subclass & gip_ins_subclass_memory_size)
                    {
                    case gip_ins_subclass_memory_word:
                    {
                        alu_mem_op = gip_mem_op_store_word;
                    }
                    case gip_ins_subclass_memory_half:
                    {
                        alu_mem_op = gip_mem_op_store_half;
                    }
                    case gip_ins_subclass_memory_byte:
                    {
                        alu_mem_op = gip_mem_op_store_byte;
                    }
                    }
                    alu_accepting_rfr_instruction_if_rfw_does = 1;
                    alu_accepting_rfr_instruction_if_mem_does = 1;
                }
                case gip_ins_class_load:
                {
                    alu_mem_rd = alu_inst.gip_ins_rd;
                    part_switch (alu_inst.gip_ins_subclass & gip_ins_subclass_memory_size)
                    {
                    case gip_ins_subclass_memory_word:
                    {
                        alu_mem_op = gip_mem_op_load_word;
                    }
                    case gip_ins_subclass_memory_half:
                    {
                        alu_mem_op = gip_mem_op_load_half;
                    }
                    case gip_ins_subclass_memory_byte:
                    {
                        alu_mem_op = gip_mem_op_load_byte;
                    }
                    }
                    alu_accepting_rfr_instruction_if_mem_does = 1;
                }
                }
            }
            else
            {
                alu_accepting_rfr_instruction_always = 1;
            }
        }

    /*b Determine pipeline results: gip_pipeline_flush, gip_pipeline_tag, gip_pipeline_executing
     */
    determine_pipeline_results "Determine pipeline results":
        {
            gip_pipeline_flush = alu_inst.f && first_cycle_of_instruction;
            gip_pipeline_executing = first_cycle_of_instruction;
            gip_pipeline_tag = alu_inst.tag;
            if (!condition_passed) // Also kills flush if the instruction is invalid
            {
                gip_pipeline_flush = 0;
                gip_pipeline_executing = 0;
            }
//            if (alu_accepting_rfr_instruction) // Also kill flush if we are blocked for actually completing the instruction - this is clearly wrong. The flush actually needs to occur as early as possible anyway.
//            {
//                gip_pipeline_flush = 0;
//                gip_pipeline_executing = 0;
//            }
        }

    /*b Copy the instruction across - alu_inst
     */
    pipeline_instruction "Pipeline instruction":
        {
            first_cycle_of_instruction <= 0;
            if (alu_accepting_rfr_instruction)
            {
                alu_inst <= rfr_inst;
                if (gip_pipeline_flush) // How do we cope with delay slots with this!!! - note that the rfr_inst may have the 'd' bit set...
                {
                    alu_inst.valid <= 0;
                }
                first_cycle_of_instruction <= 1;
            }
        }

    /*b Store flags, ALU inputs, CP indications, accumulator and shifter
     */
    alu_regs "ALU Regs":
        {
            /*b Select next values for ALU inputs based on execution blocked, or particular ALU operation (multiplies particularly)
             */
            if ( (rfr_inst.valid) &&
                 !(gip_pipeline_flush) &&
                 alu_accepting_rfr_instruction )
            {
                alu_a_in <= rf_read_port_0;
                if ( (rfr_inst.gip_ins_class==gip_ins_class_arith) &&
                     (rfr_inst.gip_ins_subclass==gip_ins_subclass_arith_mlb) )
                {
                    alu_b_in[30;2] <= alu_b_in[30;0];// An MLB instruction in RF read stage implies shift left by 2; but only if it moves to the ALU stage, which it does here
                    alu_b_in[2;0] <= 0;
                }
                elsif (rfr_inst.rm_is_imm)
                {
                    alu_b_in <= rfr_inst.immediate; // If immediate, pass immediate data in
                }
                else
                {
                    alu_b_in <= rf_read_port_1; // Else read register/special
                }
            }

            /*b Update ALU result, accumulator, shifter and flags
             */
            if ( (alu_accepting_rfr_instruction) &&
                 (alu_inst.valid) )
            {
                flags <= next_flags;
                acc <= next_acc;
                shf <= next_shf;
            }

        }

    /*b Done
     */
}
