// Pin counts
//   MII Tx 8 - TxCk, TxEn, TxD[4], TxCRS, TxCol
//   MII Rx 7 - RxCk, RxDv, RxD[4], RxEr
//  RMII Tx 6 - TxCk, TxEn, TxD[2], TxCRS, TxCol
//  RMII Rx 5 - RxCk, RxDv, RxD[2], RxEr
//  GPIO 8 - (Ck), D[8] // on receive, when an input changes it is recorded; tx is purely set/clear/write
//   SPI -
//   I2C - use GPIO
//   I2O -
//  MDIO - MDC, MDD
//HSS Tx 6 - TxCk, TxF, TxD[4] // supports T1, E1, TDM bus (1-4 bits of bus at a time), arbitrary framing inc I2S
//HSS Rx 6 - RxCk, RxF, RxD[4] // supports T1, E1, TDM bus (1-4 bits of bus at a time), arbitrary framing inc I2S
//   USB - 
//UART Tx- TxD, TxCTS, DTR
//UART Rx- RxD, RxCTS, DR
//16bD Tx 18 - TxCk, TxEn, TxD[16] // depending on mode, TxEn may be ignored, undriven or driven - bit size 1 thru 16
//16bD Rx 18 - RxCk, RxEn, RxD[16] // depending on mode, RxEn may be ignored, or driven - bit size 1 thru 16

// We want to support
// a. 2 ethernet (RMII*2)
// b. 1 ethernet (MII -  TxCk, TxEn, TxD[2], TxCrs, TxCol, RxCk, RxDv, RxD[2], RxE)

/
ethernet_tx eth0( io_clock -> eth0_tx_clock,
                    io_reset = io_reset_0,
                    data_fifo_data = tx_fifo_read_tx_data_0,
                    data_fifo_read => tx_fifo_read_toggle_0,
                    cmd_fifo_empty = tx_fifo_read_data_0,
                    cmd_fifo_data = tx_fifo_read_tx_cmd_0,
                    mii_enable => eth0_mii_enable,
                    mii_data => eth0_mii_data,
                    mii_crs = eth0_mii_crs,
                    mii_col = eth0_mii_col );
                

// implements command FIFO timers, arbitration and synch for access, buffer for tx data and cmd (32-bits each)
io_tx_arb( I/O blocks, tx_fifo_ctrl )

// 32-bit wide TX FIFO RAM, probably 2k by 32,
tx_fifo_ram (tx_fifo_ctrl, data to tx_fifo_ctrl, data in from postbus);

// takes requests from the I/O (high priority, cmd over data) and the postbus (low priority)
// and returns acknowledgements. The FIFO RAM does one access per cycle, so this is the ultimate arbiter
// Implements 4 command FIFOs and 4 data FIFOS; commands are 32+32 (time+cmd), data is 32-bit.
tx_fifo_ctrl( postbus_tx_interface, io_tx_arb )

//takes commands/data from postbus and puts in to FIFO
// also takes flow control from postbus and maps it to rx side
// also takes postbus commands from postbus target and maps to immediate FIFO status reads, FIFO resets, etc.
postbus_tx_interface( postbus_target, tx_fifo ); //  has flow control mgmt to rx side


// basically initiates transfers from FIFOs when they request it (8 events?) or when asked from tx side
postbus_rx_interface( postbus_source, rx_fifo ); // takes flow control mgmt from tx side

// takes requests from the I/O (high priority, cmd over data) and the postbus (low priority)
// and returns acknowledgements. The FIFO RAM does one access per cycle, so this is the ultimate arbiter
// Implements 4 status FIFOs and 4 data FIFOS; status is 32+32 (time+cmd) with time from this block, data is 32-bit.
rx_fifo_ctrl( postbus_tx_interface, io_tx_arb )

// 32-bit wide RX FIFO RAM, probably 2k by 32,
rx_fifo_ram (rx_fifo_ctrl, data from rx_fifo_ctrl, data out to postbus);

// implements arbitration and synch for access; note status write is 2 cycles
io_rx_arb( I/O blocks, rx_fifo_ctrl )

