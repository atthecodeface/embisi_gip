/*a Includes
 */
include "gip.h"
include "gip_internal.h"

/*a Types
 */
/*t t_reg
 */
typedef struct
{
    t_gip_word value;
} t_reg;

/*t t_rf_src
 */
typedef enum [3]
{
    rf_src_mem_result,
    rf_src_rf,
    rf_src_inst_pc,
    rf_src_alu_shf_result,
    rf_src_postbus,
    rf_src_special
} t_rf_src;

/*a Module
 */
module gip_rf( clock gip_clock,
                      input bit gip_reset,

                      input t_gip_instruction_rf dec_inst,
                      output t_gip_instruction_rf rfr_inst,

                      output bit rfr_accepting_dec_instruction_always "Asserted if the RF stage is taking a proffered instruction from the decode independent of the ALU; will be asserted if the RF stage has no valid instruction to decode currently",
                      output bit rfr_accepting_dec_instruction_if_alu_does"Asserted if the RF stage is taking a proffered instruction from the decode depending on the ALU taking the current instruction; 0 if the RF has no valid instruction, or if it has an instruction blocking on a pending register scoreboard; 1 if the RF has all the data and instruction ready for the ALU, and so depends on the ALU taking its instruction",
                      input bit rfr_accepting_dec_instruction,

                      output bit rfr_postbus_read,
                      output bit[5] rfr_postbus_read_address,
                      input t_gip_word rfr_postbus_read_data,

                      output bit rfr_special_read,
                      output bit[5] rfr_special_read_address,
                      input t_gip_word rfr_special_read_data,

                      output t_gip_word rfr_port_0,
                      output t_gip_word rfr_port_1,

                      input bit alu_inst_valid, // ALU state
                      input t_gip_ins_r alu_inst_gip_ins_rd,

                      input t_gip_ins_r alu_rd,
                      input bit alu_use_shifter,
                      input t_gip_word alu_arith_logic_result,
                      input t_gip_word alu_shifter_result,

                      input t_gip_ins_r mem_1_rd,
                      input t_gip_ins_r mem_2_rd,
                      input bit mem_read_data_valid,
                      input t_gip_word mem_read_data,

                      output bit rfw_postbus_write,
                      output bit[5] rfw_postbus_write_address,
                      output bit rfw_special_write,
                      output bit[5] rfw_special_write_address,

                      input bit gip_pipeline_flush,

                      output bit rfw_accepting_alu_rd,
                      output bit gip_pipeline_rfw_write_pc,
                      output bit[32] gip_pipeline_rfw_data
               )
{
    /*b Default clock and reset
     */
    default clock gip_clock;
    default reset gip_reset;

    /*b State in the RF read stage
     */
    clocked t_gip_instruction_rf rfr_inst_in = { valid=0,
                                              gip_ins_rn = {type=gip_ins_r_type_none, r=0},
                                              gip_ins_rd = {type=gip_ins_r_type_none, r=0},
                                              gip_ins_rm = {type=gip_ins_r_type_none, r=0},
                                              rm_is_imm = 0,
                                              k=0, a=0, f=0, d=0, pc=0, tag=0 }
                                              "Instruction in the RF read stage";

    /*b State in the RF write stage
     */
    clocked t_gip_ins_r rfw_alu_rd = { type=gip_ins_r_type_none, r=0 } "The current register to be written from an ALU path instruction";
    clocked bit         rfw_use_shifter = 0 "Asserted if alu_rd indicates a write from the shifter result not the ALU result";
    clocked t_gip_word  rfw_alu_result = 0 "Registered result of the ALU";
    clocked t_gip_word  rfw_shf_result = 0 "Registered result of the shifter";
    comb t_gip_word alu_shf_result "Mux of rfw_alu_result and rfw_shf_result, depending on rfw_use_shifter";

    clocked t_gip_ins_r rfw_mem_rd = { type=gip_ins_r_type_none, r=0 } "Type of register file write requested for the result of memory operation";
    clocked t_gip_word  rfw_mem_result = 0 "Register result of the memory stage";
    clocked bit         rfw_accepting_alu_rd = 0 "Asserted if the RFW stage can take an ALU register write; 0 only if the mem_rd is not-none and the alu_rd is not-none";

    comb t_gip_ins_r rfw_rd "Actual register being written in to the register file in this cycle";
    comb t_gip_word rfw_data "Write data being written in to the register file or other register in this cycle";

    /*b Combinatorials in the RF
     */
    comb bit rfr_blocked;
    comb bit rfw_write_enable "Asserted if the register file is to be written with the current address and data";
    comb t_rf_src read_port_0_src "Source of RF read port 0 data";
    comb t_rf_src read_port_1_src "Source of RF read port 1 data";
//    net t_gip_word rf_read_port_0 "Register file read port 0 value";
//    net t_gip_word rf_read_port_1 "Register file read port 1 value";

    /*b Instantiate register file
     */
    net bit[32] rfr_rf_data_0;
    net bit[32] rfr_rf_data_1;            
    rf_inst "":
        {

            rf_2r_1w_32_32 rf( rf_clock <- gip_clock,
                               rf_reset <= gip_reset,
                               rf_rd_addr_0 <= rfr_inst_in.gip_ins_rn.r,
                               rf_rd_data_0 => rfr_rf_data_0,
                               rf_rd_addr_1 <= rfr_inst_in.gip_ins_rm.r,
                               rf_rd_data_1 => rfr_rf_data_1,
                               rf_wr_enable <= rfw_write_enable,
                               rf_wr_addr <= rfw_rd.r,
                               rf_wr_data <= rfw_data );

            if (!rfr_inst_in.valid)
            {
                read_port_0_src = rf_src_inst_pc; // For internal results give the PC - other possibles are ACC and SHF, which will be replaced in ALU stage anyway
            }
            else
            {
                read_port_0_src = rf_src_inst_pc;
                part_switch (rfr_inst_in.gip_ins_rn.type)
                    {
                    case gip_ins_r_type_register:
                    {
                        if ( ( rfw_alu_rd.type == gip_ins_r_type_register) && (rfr_inst_in.gip_ins_rn.r == rfw_alu_rd.r ) )
                        {
                            read_port_0_src = rf_src_alu_shf_result;
                        }
                        elsif ( ( rfw_mem_rd.type == gip_ins_r_type_register) && (rfr_inst_in.gip_ins_rn.r == rfw_mem_rd.r ) )
                            {
                                read_port_0_src = rf_src_mem_result;
                            }
                        else
                        {
                            read_port_0_src = rf_src_rf;
                        }
                    }
                    case gip_ins_r_type_special:
                    {
                        read_port_0_src = rf_src_special;
                    }
                    case gip_ins_r_type_postbus:
                    {
                        read_port_0_src = rf_src_postbus;
                    }
                    }
            }

            if (!rfr_inst_in.valid)
            {
                read_port_1_src = rf_src_inst_pc; // For internal results give the PC - other possibles are ACC and SHF, which will be replaced in ALU stage anyway
            }
            else
            {
                read_port_1_src = rf_src_inst_pc;
                part_switch (rfr_inst_in.gip_ins_rm.type)
                    {
                    case gip_ins_r_type_register:
                    {
                        if ( ( rfw_alu_rd.type == gip_ins_r_type_register) && (rfr_inst_in.gip_ins_rm.r == rfw_alu_rd.r ) )
                        {
                            read_port_1_src = rf_src_alu_shf_result;
                        }
                        elsif ( ( rfw_mem_rd.type == gip_ins_r_type_register) && (rfr_inst_in.gip_ins_rm.r == rfw_mem_rd.r ) )
                            {
                                read_port_1_src = rf_src_mem_result;
                            }
                        else
                        {
                            read_port_1_src = rf_src_rf;
                        }
                    }
                    case gip_ins_r_type_special:
                    {
                        read_port_1_src = rf_src_special;
                    }
                    case gip_ins_r_type_postbus:
                    {
                        read_port_1_src = rf_src_postbus;
                    }
                    }
            }

            /*b Read the register file
             */
            rfr_port_0 = rfr_rf_data_0;
            full_switch ( read_port_0_src )
            {
            case rf_src_rf:             { rfr_port_0 = rfr_rf_data_0; }
            case rf_src_inst_pc:        { rfr_port_0 = rfr_inst_in.pc; }
            case rf_src_alu_shf_result: { rfr_port_0 = alu_shf_result; }
            case rf_src_mem_result:     { rfr_port_0 = rfw_mem_result; }
            case rf_src_postbus:        { rfr_port_0 = rfr_postbus_read_data; }
            case rf_src_special:        { rfr_port_0 = rfr_special_read_data; }
            }
            rfr_port_1 = rfr_rf_data_1;
            full_switch ( read_port_1_src )
            {
            case rf_src_rf:             { rfr_port_1 = rfr_rf_data_1; }
            case rf_src_inst_pc:        { rfr_port_1 = rfr_inst_in.pc; }
            case rf_src_alu_shf_result: { rfr_port_1 = alu_shf_result; }
            case rf_src_mem_result:     { rfr_port_1 = rfw_mem_result; }
            case rf_src_postbus:        { rfr_port_1 = rfr_postbus_read_data; }
            case rf_src_special:        { rfr_port_1 = rfr_special_read_data; }
            }
        }

    /*b Determine whether to block or not
     */
    fred "Determine whether to accept another instruction from decode":
        {
            /*b If instruction is not valid, accept instruction
             */
            rfr_accepting_dec_instruction_always = 0;
            if (!rfr_inst_in.valid)
            {
                rfr_accepting_dec_instruction_always = 1;
            }

            /*b If instruction is valid, then accept instruction only if ALU takes this and we are not blocking
             */
            rfr_blocked = 0;
            if (rfr_inst_in.valid)
            {
                if ( (rfr_inst_in.gip_ins_rn.type==gip_ins_r_type_internal) && 
                     (rfr_inst_in.gip_ins_rn.r==gip_ins_rnm_int_block_all) ) // Blocked if anything has a write pending
                {
                    if (mem_1_rd.type!=gip_ins_r_type_none)
                    {
                        rfr_blocked = 1;
                    }
                    if (mem_2_rd.type!=gip_ins_r_type_none)
                    {
                        rfr_blocked = 1;
                    }
                    if (alu_rd.type!=gip_ins_r_type_none)
                    {
                        rfr_blocked = 1;
                    }
                    if ( alu_inst_valid &&
                         (alu_inst_gip_ins_rd.type!=gip_ins_r_type_none) )
                    {
                        rfr_blocked = 1;
                    }
                }
                if (rfr_inst_in.gip_ins_rn.type==gip_ins_r_type_register) // Blocked if ALU stage will write to Rn, or memory stage will write to Rn, or our ALU holding register is for Rn
                {
                    if ( alu_inst_valid &&
                         (alu_inst_gip_ins_rd.type==gip_ins_r_type_register) &&
                         (rfr_inst_in.gip_ins_rn.r[5;0]==alu_inst_gip_ins_rd.r[5;0]) )
                    {
                        rfr_blocked = 1;
                    }
                    if ( (mem_1_rd.type==gip_ins_r_type_register) &&
                         (rfr_inst_in.gip_ins_rn.r==mem_1_rd.r) )
                    {
                        rfr_blocked = 1;
                    }
                    if ( (mem_2_rd.type==gip_ins_r_type_register) &&
                         (rfr_inst_in.gip_ins_rn.r==mem_2_rd.r) )
                    {
                        rfr_blocked = 1;
                    }
                    if ( (rfw_mem_rd.type!=gip_ins_r_type_none) &&
                         (rfw_alu_rd.type==gip_ins_r_type_register) &&
                         (rfr_inst_in.gip_ins_rn.r==rfw_alu_rd.r) )
                    {
                        rfr_blocked = 1;
                    }
                }
                if (rfr_inst_in.gip_ins_rm.type==gip_ins_r_type_register) // Blocked if ALU stage will write to Rm, or memory stage will write to Rm, or our ALU holding register is for Rm
                {
                    if ( alu_inst_valid &&
                         (alu_inst_gip_ins_rd.type==gip_ins_r_type_register) &&
                         (rfr_inst_in.gip_ins_rm.r==alu_inst_gip_ins_rd.r) )
                    {
                        rfr_blocked = 1;
                    }
                    if ( (mem_1_rd.type==gip_ins_r_type_register) &&
                         (rfr_inst_in.gip_ins_rm.r==mem_1_rd.r) )
                    {
                        rfr_blocked = 1;
                    }
                    if ( (mem_2_rd.type==gip_ins_r_type_register) &&
                         (rfr_inst_in.gip_ins_rm.r==mem_2_rd.r) )
                    {
                        rfr_blocked = 1;
                    }
                    if ( (rfw_mem_rd.type!=gip_ins_r_type_none) && // If writing something for mem stage then block if we want the ALU stage result
                         (rfw_alu_rd.type==gip_ins_r_type_register) &&
                         (rfr_inst_in.gip_ins_rm.r==rfw_alu_rd.r) )
                    {
                        rfr_blocked = 1;
                    }
                }
            }
            rfr_accepting_dec_instruction_if_alu_does = !rfr_blocked;
        }

    /*b Instruction to ALU
     */
    instruction_to_alu "Instruction to ALU":
        {
            rfr_inst = rfr_inst_in;
            rfr_inst.valid = rfr_inst_in.valid && !rfr_blocked;
        }

    /*b Postbus and special read/write
     */
    special_and_postbus "Read and write the special and postbus data":
        {
            rfr_postbus_read = 0;
            rfr_postbus_read_address = 0;
            rfr_special_read = 0;
            rfr_special_read_address = 0;
            part_switch (rfr_inst_in.gip_ins_rn.type)
                {
                case gip_ins_r_type_postbus:
                {
                    rfr_postbus_read = 1;
                    rfr_postbus_read_address = rfr_inst_in.gip_ins_rn.r;
                }
                case gip_ins_r_type_special:
                {
                    rfr_special_read = 1;
                    rfr_special_read_address = rfr_inst_in.gip_ins_rn.r;
                }
                }
            part_switch (rfr_inst_in.gip_ins_rm.type)
                {
                case gip_ins_r_type_postbus:
                {
                    rfr_postbus_read = 1;
                    rfr_postbus_read_address = rfr_postbus_read_address | rfr_inst_in.gip_ins_rm.r;
                }
                case gip_ins_r_type_special:
                {
                    rfr_special_read = 1;
                    rfr_special_read_address = rfr_special_read_address | rfr_inst_in.gip_ins_rm.r;
                }
                }
            rfw_postbus_write = 0;
            rfw_special_write = 0;
            rfw_postbus_write_address = rfw_rd.r;
            rfw_special_write_address = rfw_rd.r;
            part_switch (rfw_rd.type)
                {
                case gip_ins_r_type_special:
                {
                    rfw_special_write = 1;
                }
                case gip_ins_r_type_postbus:
                {
                    rfw_postbus_write = 1;
                }
                }
        }

    /*b Register file writeback logic - rfw_write_enable, rfw_data, rfw_read, gip_pipeline_rfw_write_pc, gip_pipeline_rfw_data
     */
    rf_writeback "Register file writeback logic":
        {
            rfw_write_enable = 0;
            if (rfw_rd.type==gip_ins_r_type_register)
            {
                rfw_write_enable = 1;
            }
            alu_shf_result = rfw_use_shifter ? rfw_shf_result : rfw_alu_result;
            rfw_data = alu_shf_result;
            rfw_rd = rfw_alu_rd;
            if (rfw_mem_rd.type!=gip_ins_r_type_none)
            {
                rfw_rd = rfw_mem_rd;
                rfw_data = rfw_mem_result;
            }

            gip_pipeline_rfw_write_pc = 0;
            if ( (rfw_rd.type==gip_ins_r_type_internal) &&
                 (rfw_rd.r==gip_ins_r_int_pc) )
            {
                gip_pipeline_rfw_write_pc = 1;
            }
            gip_pipeline_rfw_data = rfw_data;
        }

    /*b Pipeline instruction for RF read stage
     */
    pipeline_rfr_stage "Pipeline instruction for RF read stage":
        {
            if (rfr_accepting_dec_instruction)
            {
                rfr_inst_in <= dec_inst;
                if (gip_pipeline_flush)
                {
                    rfr_inst_in.valid <= 0;
                }
            }
            else // Not willing to take another instruction; we must have one on hold - flush if asked AND if it is not 'D'
            {
                if ( gip_pipeline_flush && !rfr_inst_in.d )
                {
                    rfr_inst_in.valid <= 0;
                }
            }
        }

    /*b Record RFW stage results for the write stage
     */
    pipeline_rfw_stage "Pipeline results and 'rd's for RF write stage":
        {
            if (rfw_accepting_alu_rd) // If we promised to take the next ALU rd, then take it
            {
                rfw_alu_rd <= alu_rd;
                rfw_alu_result <= alu_arith_logic_result;
                rfw_use_shifter <= alu_use_shifter;
                rfw_shf_result <= alu_shifter_result;
            }
            if (mem_read_data_valid)
            {
                rfw_mem_rd <= mem_2_rd;
                rfw_mem_result <= mem_read_data;
            }
            else
            {
                rfw_mem_rd.type <= gip_ins_r_type_none;
            }
            rfw_accepting_alu_rd <= 1;
            if ( (rfw_alu_rd.type!=gip_ins_r_type_none) ) // If we have a write to do
            {
                if ( (rfw_mem_rd.type!=gip_ins_r_type_none) ) // If we are not doing it
                {
                    rfw_accepting_alu_rd <= 0; // Then we won't be able to take another
                }
            }
        }

    /*b Done
     */
}
