/*a Includes
 */
include "gip.h"
include "gip_internal.h"
include "gip_decode.h"

/*a Types
 */
/*t t_gip_decode_state
 */
typedef fsm
{
    gip_decode_state_idle;
    gip_decode_state_native;
    gip_decode_state_emulate;
    gip_decode_state_preempt;
} t_gip_decode_state;

/*a Module
  Fetch... (for native mode... for ARM mode 'instruction blocked' should be expanded to include 'next cycle of opcode is zero')
    current instruction not valid AND prefetch not issued -> fetch current prefetch
    current instruction not valid AND prefetch issued -> fetch last prefetch
    current instruction valid AND instruction not blocked -> fetch sequential
    current instruction valid AND instruction blocked -> fetch hold
  Prefetch...
    current instruction not valid AND prefetch not issued AND pc to be valid -> prefetch new address (prefetch deemed issued)
    current instruction not valid AND prefetch issued -> prefetch sequential
    current instruction valid AND instruction blocked -> prefetch hold
    current instruction valid AND instruction not branch AND instruction not blocked -> prefetch sequential
    current instruction valid AND instruction branch AND instruction not blocked -> prefetch new address
  If flush occurs, then 'prefetch issued' is cleared in the following cycle, PC marked as invalid, and any opcode fetched is marked as invalid (prefetch deemed not issued)
  If a write of the PC occurs then the PC is to be valid; this should only occur once the prefetch is marked as not issued (after a flush)

  But... if not in native or emulate mode, then prefetch is none and fetch is hold

 */
module gip_decode( clock gip_clock,
                   input bit gip_reset,

                   output bit fetch_16,
                   output t_gip_fetch_op fetch_op, // Early in the cycle, so data may be returned combinatorially
                   input t_gip_word fetch_data,
                   input bit fetch_data_valid,
                   input bit[32] fetch_pc,
                   output t_gip_prefetch_op prefetch_op, // Late in the cycle; can be used to start an SRAM cycle in the clock edge for fetch data in next cycle (if next cycle fetch requests it)
                   output bit[32] prefetch_address,

                   output t_gip_instruction_rf dec_inst,
                   input bit rfr_accepting_dec_instruction,

                   input bit gip_pipeline_flush,
                   input bit gip_pipeline_rfw_write_pc,
                   input bit gip_pipeline_executing,
                   input bit[2] gip_pipeline_tag,
                   input t_gip_word gip_pipeline_rfw_data,

                   input bit sched_thread_to_start_valid,
                   input bit[3] sched_thread_to_start,
                   input bit[32] sched_thread_to_start_pc,
                   output bit acknowledge_scheduler,

                   input bit[8] special_repeat_count,
                   input bit[2] special_alu_mode,
                   input bit special_cp_trail_2

    )
{
    /*b Default clock and reset
     */
    default clock gip_clock;
    default reset gip_reset;

    /*b Scheduler interface
     */
    clocked bit acknowledge_scheduler=0;

    /*b Prefetch/fetch interface
     */
    clocked t_gip_word fetched_opcode = 0;
    clocked bit fetched_opcode_valid = 0;

    clocked bit valid_prefetch_issued = 0;
    clocked bit pc_valid = 0;
    clocked bit[32] pc = 0;

    /*b Decode state machine and current thread information
     */
    clocked t_gip_decode_state op_state=gip_decode_state_idle;
    clocked bit[3] thread=0;

    /*b Instruction
     */
    clocked t_gip_instruction_rf dec_inst = { valid=0,
                                              gip_ins_rn = {type=gip_ins_r_type_none, r=0},
                                              gip_ins_rd = {type=gip_ins_r_type_none, r=0},
                                              gip_ins_rm = {type=gip_ins_r_type_none, r=0},
                                              rm_is_imm = 0,
                                              k=0, a=0, f=0, d=0, pc=0, tag=0 } "Instruction in the RF read stage";
    clocked bit[5] cycle_of_opcode=0;

    /*b Accumulator tracking
     */
    clocked bit acc_valid=0;
    clocked bit[5] reg_in_acc=0;

    /*b Conditional and delay slot tracking
     */
    clocked bit in_conditional_shadow = 0;
    clocked bit in_immediate_conditional_shadow = 0;
//    clocked bit in_delay_slot = 0;
//    clocked bit follow_delay_pc = 0;
//    clocked bit[32] delay_pc=0;

    /*b Extended instruction data
     */
    clocked bit extended=0;
    clocked bit[28] extended_immediate=0;
    clocked t_gip_ins_r extended_rd={type=0,r=0};
    clocked t_gip_ins_r extended_rn={type=0,r=0};
    clocked t_gip_ins_r extended_rm={type=0,r=0};
    clocked t_gip_ext_cmd extended_cmd={extended=0};

    /*b Native instruction decoding
     */
    comb bit[16] native_opcode;
    net t_gip_instruction_rf native_dec_inst;
    net t_gip_pc_op native_dec_pc_op;
    net bit[32] native_dec_branch_offset;

    net bit native_dec_extending;
    net bit[28] native_dec_next_extended_immediate;
    net t_gip_ins_r native_dec_next_extended_rd;
    net t_gip_ins_r native_dec_next_extended_rn;
    net t_gip_ins_r native_dec_next_extended_rm;
    net t_gip_ext_cmd native_dec_next_extended_cmd;

    net bit native_dec_next_in_immediate_conditional_shadow;

    /*b Selected decode results
     */
    comb t_gip_ins_cc dec_cc;
    comb bit request_fetch;
    comb bit next_pc_valid;
    comb bit[32] next_pc;
    comb t_gip_pc_op next_pc_op;

    /*b Not implemented yet
     */
    comb bit instruction_blocked;
    comb bit branch;
    comb bit[32] branch_pc;

    /*b Not implemented
     */
    nyi "" :
        {
            instruction_blocked = 0;
            if (dec_inst.valid && !rfr_accepting_dec_instruction)
            {
                instruction_blocked = 1;
            }
            branch = 0;
            if (native_dec_pc_op==gip_pc_op_branch)
            {
                branch = 1;
            }
            branch_pc = pc + 8 + native_dec_branch_offset;
        }

    /*b Register prefetched instruction
     */
    prefetched "":
        {
            fetch_16 = 1;
            fetch_op = gip_fetch_op_this_prefetch;

            prefetch_address = next_pc;
            if (!fetched_opcode_valid)
            {
                if (!valid_prefetch_issued)
                {
                    fetch_op = gip_fetch_op_this_prefetch;
                    if (next_pc_valid)
                    {
                        prefetch_op = gip_prefetch_op_new_address;
                        prefetch_address = next_pc;
                        valid_prefetch_issued <= 1;
                    }
                    else
                    {
                        prefetch_op = gip_prefetch_op_none;
                    }
                }
                else
                {
                    fetch_op = gip_fetch_op_last_prefetch;
                    prefetch_op = gip_prefetch_op_sequential;
                }
            }
            else
            {
                if (instruction_blocked)
                {
                    fetch_op = gip_fetch_op_hold;
                    prefetch_op = gip_prefetch_op_sequential;
                }
                else
                {
                    fetch_op = gip_fetch_op_sequential; // We have an instruction decoded okay, so this is what we want; but what if the last instruction was a branch, giving new PC? We have not fetched that. Hm.
                    if (branch)
                    {
                        fetch_op = gip_fetch_op_this_prefetch; // Not if delay slot. Hmm. This is probably the issue described in the other two lines
                        prefetch_op = gip_prefetch_op_new_address;
                        prefetch_address = branch_pc;
                        valid_prefetch_issued <= 1; // So what happens in the next cycle? Instruction may not be blocked - should the fetch be 'last prefetch'?
                    }
                    else
                    {
                        prefetch_op = gip_prefetch_op_sequential;
                    }
                }
            }
            // If the prefetch_op is sequential then we can speculate a fetch also
            if (gip_pipeline_flush)
            {
                valid_prefetch_issued <= 0;
                prefetch_op = gip_prefetch_op_none;
            }

            if (!fetched_opcode_valid || !instruction_blocked)
            {
                fetched_opcode <= fetch_data;
                fetched_opcode_valid <= fetch_data_valid;
                pc <= fetch_pc;
            }
        }

    /*b Native decode - use top or bottom half of instruction (pc bit 1 is set AND native AND valid)
     */
    native_decode "":
        {
            dec_cc = gip_ins_cc_always;
            if (in_conditional_shadow)
            {
                dec_cc = gip_ins_cc_cp;
            }
            native_opcode = fetched_opcode[16;0];
            if ( (op_state!=gip_decode_state_native) || (!pc[1]) )
            {
                native_opcode = fetched_opcode[16;0];
            }
            else
            {
                native_opcode = fetched_opcode[16;16];
            }
            gip_decode_native native( opcode <= native_opcode,

                                      dec_cc <= gip_ins_cc_always, // If in ARM mode should use its condition

                                      special_repeat_count <= special_repeat_count,
                                      special_alu_mode <= special_alu_mode,

                                      inst => native_dec_inst,
                                      pc_op => native_dec_pc_op,
                                      native_mapped_branch_offset => native_dec_branch_offset,

                                      extended <= extended,
                                      extended_immediate <= extended_immediate,
                                      extended_rd <= extended_rd,
                                      extended_rn <= extended_rn,
                                      extended_rm <= extended_rm,
                                      extended_cmd <= extended_cmd,

                                      extending => native_dec_extending,
                                      next_extended_immediate => native_dec_next_extended_immediate,
                                      next_extended_rd => native_dec_next_extended_rd,
                                      next_extended_rn => native_dec_next_extended_rn,
                                      next_extended_rm => native_dec_next_extended_rm,
                                      next_extended_cmd => native_dec_next_extended_cmd,

                                      in_conditional_shadow <= in_conditional_shadow,
                                      in_immediate_conditional_shadow <= in_immediate_conditional_shadow,
                                      next_in_immediate_conditional_shadow => native_dec_next_in_immediate_conditional_shadow );
        }

    /*b Handle according to operating state
     */
    decode_state_machine "Handle according to operating state":
        {
            dec_inst <= native_dec_inst;
            request_fetch = 0;
            next_pc_valid = 0;
            next_pc = 0;
            acknowledge_scheduler <= 0;
            full_switch (op_state)
            {
                /*b Idle - wait for schedule request
                 */
            case gip_decode_state_idle:
            {
                if (sched_thread_to_start_valid)
                {
                    op_state <= gip_decode_state_native;
                    acknowledge_scheduler <= 1;
                    thread <= sched_thread_to_start;
                    next_pc = sched_thread_to_start_pc;
                    next_pc_valid = 1;
                }
                acc_valid <= 0;
                cycle_of_opcode <= 0;
                in_conditional_shadow <= 0;
                in_immediate_conditional_shadow <= 0;
                extended_immediate <= 0;
                extended_cmd.extended <= 0;
                extended_rd.type <= gip_ins_r_type_no_override;
                extended_rn.type <= gip_ins_r_type_no_override;
                extended_rm.type <= gip_ins_r_type_no_override;
                dec_inst.valid <= 0;
            }
            /*b Native - decode top or bottom half of instruction (pc bit 1 is set AND native AND valid)
             */
            case gip_decode_state_native:
            {
                /*b Select native instruction as our decode
                 */
                if (rfr_accepting_dec_instruction)
                {
                    dec_inst <= native_dec_inst;
                    dec_inst.pc <= pc;
                    if (!fetched_opcode_valid)
                    {
                        dec_inst.valid <= 0;
                    }
                    else
                    {
                        next_pc_op = native_dec_pc_op;
                        cycle_of_opcode <= 0;

//                    acc_valid <= next_acc_valid;
//                    reg_in_acc <= next_reg_in_acc;

                        extended_immediate <= native_dec_next_extended_immediate;
                        extended_cmd <= native_dec_next_extended_cmd;
                        extended_rd <= native_dec_next_extended_rd;
                        extended_rn <= native_dec_next_extended_rn;
                        extended_rm <= native_dec_next_extended_rm;

                        in_conditional_shadow <= 0;
                        in_immediate_conditional_shadow <= 0;
                        if (native_dec_next_in_immediate_conditional_shadow)
                        {
                            in_conditional_shadow <= 1;
                            in_immediate_conditional_shadow <= 1;
                        }
                        if ( (in_immediate_conditional_shadow) && (special_cp_trail_2) )
                        {
                            in_conditional_shadow <= 1;
                        }

//                        if (follow_delay_pc)
//                        {
//                            next_pc = delay_pc;
//                        }
                        if (!native_dec_extending)
                        {
                            extended_immediate <= 0;
                            extended_cmd.extended <= 0;
                            extended_rd.type <= gip_ins_r_type_no_override;
                            extended_rn.type <= gip_ins_r_type_no_override;
                            extended_rm.type <= gip_ins_r_type_no_override;
                        }

                        if (gip_pipeline_rfw_write_pc)
                        {
                            next_pc = gip_pipeline_rfw_data;
                            next_pc_valid = 1;
                        }
                        if (gip_pipeline_flush)
                        {
                            pc_valid <= 0;
                            acc_valid <= 0;

                            extended_immediate <= 0;
                            extended_cmd.extended <= 0;
                            extended_rd.type <= gip_ins_r_type_no_override;
                            extended_rn.type <= gip_ins_r_type_no_override;
                            extended_rm.type <= gip_ins_r_type_no_override;

                            dec_inst.valid <= 0;
//                            in_delay_slot <= 0;
//                            follow_delay_pc <= 0;
                            in_immediate_conditional_shadow <= 0;
                            in_conditional_shadow <= 0;
                        }
                        if (gip_pipeline_tag && gip_pipeline_executing)
                        {
                            op_state <= gip_decode_state_idle;
                        }
                    }
                }
            /*b All done
             */
            }
        }
    }
}

