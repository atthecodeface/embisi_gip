/*a Includes
 */
include "gip.h"
include "gip_internal.h"

/*a Types
 */

/*a Module
 */
module gip_alu_barrel_shift( input bit carry_in,
                             input t_gip_shift_op gip_shift_op,
                             input t_gip_word value,
                             input bit[8] amount,
                             output t_gip_word result,
                             output bit carry_out )
    "
This module implements a 5-operation barrel shifter.

It takes a 32-bit data input with carry, performs a shift or rotate,
and produces a 32-bit result with carry out.

The amount of the shift is a value from 0 to 255; a shift of 0 is deemed
to be no shift at all, and the carry out is the same as the carry in.

Now, imagine we are shifting not a 32-bit number, but a 4-bit number 'abcd'

We are going to implement the shifter with a 4-bit barrel shift. We also generate a mask dependent on the amount

Amt / -amt   BR       Mask
  0 / 4     abcd     1111
  1 / 3     dabc     0111
  2 / 2     cdab     0011
  3 / 1     bcda     0001
  4 / 0     abcd     0000

LSL(-amt) is BR & ~Mask, with carry BR[0]
LSR(amt)  is BR & Mask, with carry BR[3]
ASR(amt)  is a?BR|~Mask:BR&Mask, with carry BR[3]
ROR(amt)  is BR, with carry BR[3]
RRX       is Cin.BR[3;0], with carry BR[0]

Note that RRX is called with amount==32 for ARM instructions

"
{
    comb bit[8] rot_amount;
    comb t_gip_word value_rot_stage_1;
    comb t_gip_word value_rot_stage_2;
    comb t_gip_word value_rot_stage_3;
    comb t_gip_word value_rot_stage_4;
    comb t_gip_word value_rot_stage_5;
    comb t_gip_word barrel_shift_result;
    comb t_gip_word mask;
    comb bit[4] mask_bottom_bits;

    /*b rot_amount
     */
    rot_amount "Calculate rotate amount":
        {
            // ror(0) gives mask ffff
            // ror(1) gives mask 7fff
            // ror(31) gives mask 1
            // ror(32) gives mask 0
            // ror(>32) gives mask 0
            rot_amount = amount;
            if (gip_shift_op==gip_shift_op_lsl)
            {
                // want... 
                // lsl(0)=>ror(32),mask=0     => same as ror(32)
                // lsl(1)=>ror(31),mask=1     => same as ror(31)
                // lsl(31)=>ror(1),mask=7fff  => same as ror(1)
                // lsl(32)=>ror(0),mask=ffff  => same as ror(0)
                // lsl(>32)=>ror(x),mask=x (picked up as a special case later)
                rot_amount = 32-amount;
            }
            if (gip_shift_op==gip_shift_op_rrx) // ensure rrx is rotate by 1, as amount in should be 32
            {
                rot_amount[0] = 1;
            }
        }

    /*b Barrel shift and mask
     */
    barrel_shift_and_mask "Barrel shifter and mask generation":
        {
            /*b Mask - set bottom (31-rot_amount) bits, or rather clear top rot_amount bits
             */
            full_switch(rot_amount[2;0])
            {
            case 0: {mask_bottom_bits = 4b1111;}
            case 1: {mask_bottom_bits = 4b0111;}
            case 2: {mask_bottom_bits = 4b0011;}
            case 3: {mask_bottom_bits = 4b0001;}
            }
            full_switch(rot_amount[3;2])
            {
            case 0: {mask = 32h0fffffff; mask[4;28]=mask_bottom_bits; }
            case 1: {mask = 32h00ffffff; mask[4;24]=mask_bottom_bits; }
            case 2: {mask = 32h000fffff; mask[4;20]=mask_bottom_bits; }
            case 3: {mask = 32h0000ffff; mask[4;16]=mask_bottom_bits; }
            case 4: {mask = 32h00000fff; mask[4;12]=mask_bottom_bits; }
            case 5: {mask = 32h000000ff; mask[4; 8]=mask_bottom_bits; }
            case 6: {mask = 32h0000000f; mask[4; 4]=mask_bottom_bits; }
            case 7: {mask = 32h00000000; mask[4; 0]=mask_bottom_bits; }
            }
            if (rot_amount[3;5])
            {
                mask=0;
            }

            /*b Barrel shift
             */
            value_rot_stage_1 = value;
            if (rot_amount[4])
            {
                value_rot_stage_1[16; 0] = value[16;16];
                value_rot_stage_1[16;16] = value[16; 0];
            }
            value_rot_stage_2 = value_rot_stage_1;
            if (rot_amount[3])
            {
                value_rot_stage_2[24; 0] = value_rot_stage_1[24; 8];
                value_rot_stage_2[ 8;24] = value_rot_stage_1[ 8; 0];
            }
            value_rot_stage_3 = value_rot_stage_2;
            if (rot_amount[2])
            {
                value_rot_stage_3[28; 0] = value_rot_stage_2[28; 4];
                value_rot_stage_3[ 4;28] = value_rot_stage_2[ 4; 0];
            }
            value_rot_stage_4 = value_rot_stage_3;
            if (rot_amount[1])
            {
                value_rot_stage_4[30; 0] = value_rot_stage_3[30; 2];
                value_rot_stage_4[ 2;30] = value_rot_stage_3[ 2; 0];
            }
            value_rot_stage_5 = value_rot_stage_4;
            if (rot_amount[0])
            {
                value_rot_stage_5[31; 0] = value_rot_stage_4[31; 1];
                value_rot_stage_5[ 1;31] = value_rot_stage_4[ 1; 0];
            }
            barrel_shift_result = value_rot_stage_5;
        }

    /*b result and carry out
     */
    result_and_carry_out "Result and carry out determination":
        {
            result = barrel_shift_result;
            carry_out = barrel_shift_result[31];
            full_switch (gip_shift_op)
            {
            case gip_shift_op_lsl:
            {
                result = barrel_shift_result & ~mask;
                carry_out = barrel_shift_result[0];
            }
            case gip_shift_op_lsr:
            {
                result = barrel_shift_result & mask;
                carry_out = barrel_shift_result[31];
            }
            case gip_shift_op_asr:
            {
                result = value[31] ? (barrel_shift_result | ~mask) : (barrel_shift_result & mask);
                carry_out = barrel_shift_result[31];
            }
            case gip_shift_op_ror:
            {
                result = barrel_shift_result;
                carry_out = barrel_shift_result[31];
            }
            case gip_shift_op_rrx:
            {
                result = barrel_shift_result;
                result[31] = carry_in;
                carry_out = barrel_shift_result[31];
            }
            }
            if (amount==32) // ror,rrx normal; lsl=0 (already, as rot_amt==0, mask=1s); lsr=0 (already, as mask=0s); asr=all top bit (already, as mask=0s)
            {
                result=result;
            }
            elsif (amount==0) // ALWAYS PASS C and value through untouched
            {
                result = value;
                carry_out = carry_in;
            }
            elsif (amount[3;5]!=0) // 33 to 255 - override carry for lsl, lsr, asr; ror and rrx are already okay
                {
                    part_switch (gip_shift_op)
                        {
                        case gip_shift_op_lsl: {carry_out = 0; result=0;}
                        case gip_shift_op_lsr: {carry_out = 0; result=0;}
                        case gip_shift_op_asr: {carry_out = value[31]; result=value[31]?32hffffffff:0;}
                        }
                }
        }
}
