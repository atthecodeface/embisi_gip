
module utopia_pos_tx_fsm(
	clock port_clock,
	input bit port_reset,
	input bit io_cmd_fifo_ne,
	input bit io_cmd_inc_hec,
	input bit io_cmd_num_bytes,
	input bit io_cmd_drive_en_all_cell,
	input bit device_cl_av,
	input bit grant_tx_address_ctl,
	output bit io_cmd_toggle,
	output bit io_cmd_type,
	output bit next_utopia_tx_en,
	output bit next_utopia_tx_soc,
	output bit next_utopia_tx_eop,
	output bit next_utopia_td_src,
	output bit request_tx_addr_ctl 
	)
"This module supports SPHY and MPHY master Utopia TX and SPI-3 8-bit SPHY/MPHY TX, with the actual polling supported in a companion module - this module will send a cell to the given PHY using a cell available handshakepresenting the requested PHY number, but during transmission it expects someone else to do the polling of availability of other PHYs."
{
	default clock port_clock;
	default reset port_reset;
	clocked bit io_cmd_toggle=0;
	clocked bit io_cmd_type = 0;
	clocked t_utopia_tx_fsm_state fsm_state=idle;
	comb utopia_tx_fsm_state next_fsm_state;
	comb bit toggle_io_cmd;

	toggle_io_cmd = 0;
	next_fsm_state = fsm_state;
	next_utopia_tx_en = 0;
	next_utopia_tx_soc = 0;
	next_utopia_tx_eop = 0;
	switch fsm_state
	{
	case idle:
		if (io_cmd_fifo_ne)
		{
			next_fsm_state = eading_cmd_1;
			toggle_io_cmd = 1;
		}
		break;
	case reading_cmd_1:
		next_fsm_state = requesting_tx_address;
		break;
	case requesting_tx_address:
		if (grant_tx_address_ctl)
		{
			next_fsm_state = driving_address_with_data_coming;
			toggle_io_cmd = 1;
		}
		break;
	case driving_address_with_data_coming:
		if (device_cl_av)
		{
			next_fsm_state = prestart_cell;
		}
		else
		{
			next_fsm_state = drive_address_with_data_ready;
		}
		break;
	case drive_address_with_data_ready:
		next_fsm_state = driving_address_with_data_ready;
		break;
	case driving_address_with_data_ready:
		if (device_cl_av)
		{
			next_fsm_state = prestart_cell;
		}
		else
		{
			next_fsm_state = drive_address_with_data_ready;
		}
		break;
	case prestart_cell:
		berak;
	}

	if (toggle_io_cmd)
	{
		io_cmd_toggle <= !io_cmd_toggle;
	}
}



