constant integer baud_divider_size=15;

module baud_rate_generator( clock io_clock,
                            input bit io_reset,
                            output bit baud_clock_enable,
                            input bit set_clock_config,
                            input bit[baud_divider_size] config_baud_addition_value,
                            input bit[baud_divider_size] config_baud_subtraction_value )
"This is a simple-ish baud rate generator that utilizes
an error function to generate a baud clock enable.
It contains a current 'error' value that, on every clock tick,
is either:
 reduced by a number (the subtraction constant)
 or increased by a different number (the addition constant)
The sign of the 'error' value determines which of the two is performed.
If the 'error' value is negative then the addition constant is used, in an
attempt to get the 'error' value back to zero.
If the 'error' value is positive then the subtraction constant is used.
As a result, the 'error' value will oscillate around zero, spending
a certain amount of its time negative, and a certain amount positive,
with an even distribution.
The baud_clock_enable signal is asserted if the 'error' value
is non-negative.
When the addition and subtraction values are written, the
error value is also written, to the value in the subtraction constant.
To reduce gate count there is in fact only a single adder, and the
subtraction constant presented should actually be a two's complement
of the value to subtract (this save two's complement logic in hardware).

Note:
The %age of the time that the error value is nonnegative is (addc)/(subc+addc)*100.
For example, if the subtraction constant (suc) is 3, and the addition constant is 5, then
the error value runs through the following sequence:
-3 2 -1 4 1 -2 3 0   -3 2 -1 4 1 -2 3 0 ...
This is nonnegative for 5 of every 8 cycles, or (5)/(3+5)

To configure the baud enable as a simple clock divider, the addition constant should be 1
and the subtraction constant should be one less than the divider required. For example, divide by 10
with subc=9, addc=1:
-9 -8 -7 -6 -5 -4 -3 -2 -1 0   -9 -8 -7 -6 -5 -4 -3 -2 -1 0 ...

For divide by 3.3333 (or 10/3) we need subc+addc=10, addc=3 => subc=7:
-7 -4 -1 2 -8 -5 -2 1 -6 -3 0   -7 -4 -1 2 -8 -5 -2 1 -6 -3 0  ...
producing a non negative number after 4, 3, 3 4, 3, 3, 4, 3, 3... cycles,
for and average of 3.333

The error value needs to be able to divide 200MHz down to 16*1200 for 1200 baud UARTs,
so we need to be able to divide by up to 2e8/1.6e1/1.2e3 = 1.1e4 (or thereabouts) = 11,000
This implies at least 14 bits of magnitude.
For such a divider try subc=0x2af7, addc=1.
Because we need the two's complement of subc, we have two options: use an additional
magnitude bit in the error value and the constants to support the sign, or just extend the
error value for the sign and assume the top bit of the addition constant will be zero and the
top bit of the subtraction constant will be 1.

Now we have two additional requirements: a constant 'on' baud enable and a constant 'off' baud
enable. The second can be achieved with a non-zero subtraction constant and a zero addition
constant - then the error value will hold a negative value. The first can be achieved if the
subtraction constant is zero and the addition constant is zero.

With this additional constraint it is clear that we need to expand the subtraction constant
and the error value; we will also extend the addition constant for symmetry and ease-of-comprehension.

So, we need to support +-11,000 in the error value and the constants, so 15 bits of each (+-16384).
"
{
     default clock io_clock;
     default reset io_reset;

     clocked bit[baud_divider_size] baud_addition_value = 0;
     clocked bit[baud_divider_size] baud_subtraction_value = 0;
     clocked bit[baud_divider_size] baud_error_value = 0;
     clocked bit baud_clock_enable = 0;

     comb bit[baud_divider_size] baud_error_value_adder_input "Selected value of either addition or subtraction constant";
     comb bit[baud_divider_size] next_baud_error_value "Result of error function algorithm";

     configure_clock "Write the clock configuration":
          if (set_clock_config)
          {
               baud_addition_value <= config_baud_addition_value;
               baud_subtraction_value <= config_baud_subtraction_value;
          }

     next_error_value "Next error value, normal running":
          baud_error_value_adder_input = config_baud_subtraction_value;
          if (baud_error_value[baud_divider_size-1])
          {
               baud_error_value_adder_input = config_baud_addition_value;
          }
          next_baud_error_value = baud_error_value + baud_error_value_adder_input;

     counter "Baud counter and enable":
          if (set_clock_config)
          {
               baud_error_value <= config_baud_addition_value;
               baud_clock_enable <= ~config_baud_addition_value[baud_divider_size-1];
          }
          else
          {
               baud_error_value <= next_baud_error_value;
               baud_clock_enable <= next_baud_error_value[baud_divider_size-1];
          }
}
