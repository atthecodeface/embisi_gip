/*a Includes
 */
include "gip.h"
include "gip_internal.h"

/*a Types
 */

/*a Submodules
 */
/*m gip_alu_barrel_shift_data_path
 */
extern module gip_alu_barrel_shift_data_path( clock gip_clock,
                                              input bit gip_reset,
                                              input t_gip_word value,
                                              input bit[5] rotate_amount,
                                              input bit zero_mask, // if 1, zero the mask, else use top 'rotate_amount' bits of 0
                                              input bit negate_mask, // if 1,
                                              input bit and_mask, // if 0, OR the (negated) (zeroed) mask
                                              output t_gip_word result,
                                              output bit barrel_shift_bit_31,
                                              output bit barrel_shift_bit_0 )
{
    timing comb input value, rotate_amount, zero_mask, negate_mask, and_mask;
    timing comb output result, barrel_shift_bit_31, barrel_shift_bit_0;
}


/*a Module
 */
module gip_alu_barrel_shift( clock gip_clock,
                             input bit gip_reset,
                             input bit carry_in,
                             input t_gip_shift_op gip_shift_op,
                             input t_gip_word value,
                             input bit[8] amount,
                             output t_gip_word result,
                             output bit carry_out )
    "
This module implements a 5-operation barrel shifter.

It takes a 32-bit data input with carry, performs a shift or rotate,
and produces a 32-bit result with carry out.

The amount of the shift is a value from 0 to 255; a shift of 0 is deemed
to be no shift at all, and the carry out is the same as the carry in.

Now, imagine we are shifting not a 32-bit number, but a 4-bit number 'abcd'

We are going to implement the shifter with a 4-bit barrel shift. We also generate a mask dependent on the amount

Amt / -amt   BR       Mask
  0 / 4     abcd     1111
  1 / 3     dabc     0111
  2 / 2     cdab     0011
  3 / 1     bcda     0001
  4 / 0     abcd     0000

LSL(-amt) is BR & ~Mask, with carry BR[0]
LSR(amt)  is BR & Mask, with carry BR[3]
ASR(amt)  is a?BR|~Mask:BR&Mask, with carry BR[3]
ROR(amt)  is BR, with carry BR[3]
RRX       is Cin.BR[3;0], with carry BR[0]

Note that RRX is called with amount==32 for ARM instructions

"
{
    comb bit[8] rot_amount;

    comb bit zero_mask; // if 1, zero the mask, else use top 'rotate_amount' bits of 0
    comb bit negate_mask; // if 1,
    comb bit and_mask; // if 0, OR the (negated) (zeroed) mask
    net t_gip_word masked_barrel_shift;
    net bit barrel_shift_bit_31;
    net bit barrel_shift_bit_0;

    /*b rot_amount
     */
    rot_amount "Calculate rotate amount":
        {
            // ror(0) gives mask ffff
            // ror(1) gives mask 7fff
            // ror(31) gives mask 1
            // ror(32) gives mask 0
            // ror(>32) gives mask 0
            rot_amount = amount;
            if (gip_shift_op==gip_shift_op_lsl)
            {
                // want... 
                // lsl(0)=>ror(32),mask=0     => same as ror(32)
                // lsl(1)=>ror(31),mask=1     => same as ror(31)
                // lsl(31)=>ror(1),mask=7fff  => same as ror(1)
                // lsl(32)=>ror(0),mask=ffff  => same as ror(0)
                // lsl(>32)=>ror(x),mask=x (picked up as a special case later)
                rot_amount = 32-amount;
            }
            if (gip_shift_op==gip_shift_op_rrx) // ensure rrx is rotate by 1, as amount in should be 32
            {
                rot_amount[0] = 1;
            }
        }

    /*b data path controls
     */
    data_path_control "Data path controls":
        {
            /*b Defaults for ROR
             */
            zero_mask = 1;
            negate_mask = 0;
            and_mask = 0;

            /*b Choose based on op
             */
            full_switch (gip_shift_op)
            {
            case gip_shift_op_lsl: // output = barrel & ~mask
            {
                zero_mask = 0;
                negate_mask = 1;
                and_mask = 1;
                if (amount==0) // == 0, LSL is barrel & ~0
                {
                    zero_mask = 1;
                    negate_mask = 1;
                    and_mask = 1;
                }
                if (amount[3;5]!=0) // >= 32, LSL is zero = barrel & 0
                {
                    zero_mask = 1;
                    negate_mask = 0;
                    and_mask = 1;
                }
            }
            case gip_shift_op_lsr:
            {
                zero_mask = 0;
                negate_mask = 0;
                and_mask = 1;
                if (amount==0) // == 0, LSR is barrel & ~0
                {
                    zero_mask = 1;
                    negate_mask = 1;
                    and_mask = 1;
                }
                if (amount[3;5]!=0) // >= 32, LSR is zero = barrel & 0
                {
                    zero_mask = 1;
                    negate_mask = 0;
                    and_mask = 1;
                }
            }
            case gip_shift_op_asr:
            {
                if (value[31]==0) // ASR of +ve is same as LSR
                {
                    zero_mask = 0;
                    negate_mask = 0;
                    and_mask = 1;
                    if (amount==0) // == 0, ASR is barrel & ~0
                    {
                        zero_mask = 1;
                        negate_mask = 1;
                        and_mask = 1;
                    }
                    if (amount[3;5]!=0) // >= 32, ASR of +ve is zero = barrel & 0
                    {
                        zero_mask = 1;
                        negate_mask = 0;
                        and_mask = 1;
                    }
                }
                else // ASR of -ve is barrel | ~mask
                {
                    zero_mask = 0;
                    negate_mask = 1;
                    and_mask = 0;
                    if (amount==0) // == 0, ASR is barrel & ~0
                    {
                        zero_mask = 1;
                        negate_mask = 1;
                        and_mask = 1;
                    }
                    if (amount[3;5]!=0) // >= 32, ASR -ve is all 1s = barrel | 1
                    {
                        zero_mask = 1;
                        negate_mask = 1;
                        and_mask = 0;
                    }
                }
            }
            case gip_shift_op_ror:
            {
                // use barrel | 0
                zero_mask = 1;
                negate_mask = 0;
                and_mask = 0;
            }
            case gip_shift_op_rrx:
            {
                // use barrel | 0
                zero_mask = 1;
                negate_mask = 0;
                and_mask = 0;
            }
            }
        }

    /*b Data path
     */
    data_path "Data path instantiation":
        {
            gip_alu_barrel_shift_data_path data_path( gip_clock <- gip_clock,
                                                      gip_reset <= gip_reset,
                                                      value <= value,
                                                      rotate_amount <= rot_amount[5;0],
                                                      zero_mask <= zero_mask,
                                                      negate_mask <= negate_mask,
                                                      and_mask <= and_mask,
                                                      result => masked_barrel_shift,
                                                      barrel_shift_bit_31 => barrel_shift_bit_31,
                                                      barrel_shift_bit_0 => barrel_shift_bit_0 );
        }

    /*b result and carry out
     */
    result_and_carry_out "Result and carry out determination":
        {
            result = masked_barrel_shift;
            carry_out = barrel_shift_bit_31;
            part_switch (gip_shift_op)
            {
            case gip_shift_op_lsl:
            {
                carry_out = barrel_shift_bit_0;
            }
            case gip_shift_op_rrx:
            {
                result[31] = carry_in;
            }
            }
            if (amount==0) // ALWAYS PASS C and value through untouched
            {
                carry_out = carry_in;
            }
            if ((amount[3;5]!=0) && (amount!=32))
            {
                part_switch (gip_shift_op)
                {
                case gip_shift_op_lsl:
                case gip_shift_op_lsr:
                {
                    carry_out = 0;
                }
                case gip_shift_op_asr:
                {
                    carry_out = value[31];
                }
                }
            }
        }
}
