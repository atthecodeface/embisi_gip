/*a Copyright Gavin J Stark, 2004
 */

/*a To do
  Add collision handling? This is handled with mii_err
 */

/*a Includes
 */
include "io_cmd.h"
include "io_ethernet_rx.h"

/*a Constants
 */

/*a Types
 */
/*t t_data_fsm
 */
typedef fsm {
    data_fsm_idle "Idle data state, waiting for receive data";
    data_fsm_wait_for_end_of_sfd               "Waiting for end of SFD; the count indication will reach 2 when the SFD completes";
    data_fsm_reading_data                      "Reading data, calculating FCS;";
    data_fsm_reading_data_last_nybble_of_word  "Reading data, calculating FCS, write data to FIFO, possibly write status";
    data_fsm_packet_complete_waiting           "Packet complete, checked FCS, waiting for any previous data and status to have been written";
    data_fsm_packet_complete                   "Packet complete, writing final data and status";
    data_fsm_framing_error                     "Framing error (error received, data valid went away unexpectedly, etc)";
} t_data_fsm;

/*t t_data_fsm_data
 */
typedef struct 
{
    t_data_fsm state;
    bit[3] counter;
    bit[6] bytes_in_block;
    bit[10] blocks_in_packet;
} t_data_fsm_data;

/*t t_status_to_write
 */
typedef enum [3]
{
    status_to_write_block,
    status_to_write_packet_fcs_ok,
    status_to_write_packet_fcs_bad,
    status_to_write_fifo_overrun,
    status_to_write_odd_nybbles,
    status_to_write_rx_err,
    status_to_write_etx_passthrough
} t_status_to_write;

/*t t_sync
 */
typedef struct
{
    bit metastable;
    bit stable;
    bit last;
} t_sync;

/*a io_ethernet_rx module
 */
module io_ethernet_rx( clock io_clock,
                       input bit io_reset,

                       output bit[32] data_fifo_data,
                       output bit data_fifo_toggle,
                       input bit data_fifo_full,

                       output bit[32] status_fifo_data,
                       output bit status_fifo_toggle,

                       input bit mii_dv, // goes high during the preamble OR at the latest at the start of the SFD
                       input bit mii_err, // if goes high with dv, then abort the receive; wait until dv goes low
                       input bit[4] mii_data,

                       input bit etx_status_fifo_toggle, // for passing etx status through to our fifo
                       input bit[32] etx_status_fifo_data,

                       input bit[2] cfg_padding
 )

    /*b Documentation
     */
"
This module implements an I/O target to ethernet MII/RMII receive conversion. It utilizes a single status FIFO to indicate if received packets have an even number of nybbles, if the CRC is correct, and if the framing is correct (SFD, no errors in packet). Data is put in to the data FIFO 32-bits at a time. Every 64 bytes a status is presented, indicating that the packet is complete or there should be more to come.

The receive inputs are registered on entry to the system.

The basic structure is a single state machine, with a counter that counts the residence time in that state.
It starts off idle, and when data is received the state machine checks for preamble, then SFD (exactly 2 nybbles); it then pumps data in to a 32-bit storage register which is pushed to the data FIFO, counting the bytes. When the 64th byte is being pushed in a status word is also sent. When the end of the packet is reached a further status is sent indicating the size of the last block.

This flow means that every nybble from just after the SFD to the final nybble of the FCS is sent. The FCS valid indication is included in the final status of a packet

FIFO OVERRUN? Do not let the FIFO overrun, as the best approach; however, data fifo overrun is indicated in the status, and is detected if we issue a write to the data FIFO when it indicates full: note that this means protecting the status FIFO from overrun is most important if any overrun can occur

1. Idle
2. valid data received (without error), preamble or sfd -> wait for end of sfd; if data valid and error, or data valid and not preamble or sfd indication, then it is a framing error
3. wait for end of sfd
4. store nybbles, calculate FCS, until 7 nybbles received; then go to 5. However, if not data valid, go to state 6 (if even nybbles received) or framing error (if odd nybbles received)
5. store eighth nybble, calculate FCS; copy to storage register, increment words written, and write to data FIFO; if 16 words written write status also; go back to 4. However, if not data valid then hit framing error instead (as half-way through a byte)

6. Wanted to store an odd nybble in the holding register, but it was not valid; must be end of packet! Record 'FCS correct' status. Record length of packet. Wait in this state for up to 8 counts, shifting data up (also for last status and data to be written).
7. Send final word of data to FIFO (if there is some), and write status; wait for 8 clocks, then return to idle.

Framing errors occurring in the packet or data FIFO overun (bad SFD, data valid going away mid-byte) cause the framing error state to be entered; this sends a status message indicating the number of words written, and the reason for the framing error; it waits for 8 cycles then returns to idle.


The status from the etx can be piped in through here to allow a full ethernet to run on a single IO slot
To do this the etx status must be written when the rx will not require the bus
Now, the rx will only write a status for completion or error after sitting in the data_fsm_packet_complete or data_fsm_framing_error states for 8 clocks, so we do not pass through in those states
Also the rx may write out a block complete if it is in data_fsm_reading_data or data_fsm_reading_data_last_nybble_of_word and the bytes in the block indicates block completion, so we must avoid that.
So we pass through etx in the following circumstances:
 idle and its been >8 ticks since status (to allow for other status to be written)
 wait_for_end_of_sfd and its been >8 cycles since status
 data (inc last nybble of word) and its been >8 ticks since status and we are >8 ticks (nybbles) = 4 bytes before the end of a block (bytes_in_block<60)

"
{

    /*b Clock and reset
     */
    default clock io_clock;
    default reset io_reset;

    /*b MII registers
     */
    clocked bit[4] r_mii_rx_data = 0;
    clocked bit    r_mii_rx_dv = 0;
    clocked bit    r_mii_rx_err = 0;

    /*b State and combinatorials for the data FSM
     */
    clocked   t_data_fsm_data   data_fsm = {state=data_fsm_idle, counter=0, bytes_in_block=0, blocks_in_packet=0} "Actual FSM state the receive data FSM is in";
    comb   t_data_fsm_data      next_data_fsm "Next state for the data FSM";
    comb bit word_complete      "Indicates a word needs to be written to the data FSM";

    /*b State and combinatorials for the data path, including FCS
     */
    comb      bit[4]        data_for_fcs "Data nybble XOR FCS bits that are the effective feedback into the FCS calculation";
    clocked   bit[32]       fcs = 32hffffffff "FCS store, initialized to all 1's";
    comb      bit[32]       next_fcs "Combinatorial value for next FCS, particularly during calculation: may be overridden by initialization or shift-register values";
    comb      bit           fcs_ok "Asserted if the current FCS value indicates a correct FCS for a packet";

    clocked bit[32] data_register = 0;
    comb bit[32] next_data_register;
    clocked bit[32] data_fifo_data = 0 "Data to write to the data fifo";
    clocked bit data_fifo_toggle = 0 "Toggled to indicate that the data in data_fifo_data should be written to the data FIFO";

//    clocked bit[32] status_fifo_data = 0 "Data to write to status FIFO";
    clocked bit status_fifo_toggle = 0 "Toggled to indicate a write to the status FIFO should occur";
    clocked bit status_write = 0 "Asserted if we should write status to the status FIFO; should always have at least 7 clock ticks between assertions";
    clocked t_status_to_write status_to_write = status_to_write_block      "Status we should write if status_write is high";
    clocked t_status_to_write status_being_written = status_to_write_block "Status type we are writing";
    clocked bit[3]status_wait = 0 "If non-zero then must wait before writing status (for etx particularly - the rest should be clean by design)";

    comb bit status_block_etx_passthrough "Asserted if etx status data cannot be written as other status has been or may be";
    comb bit status_write_passthrough "Asserted if etx status data should be written";
    clocked bit status_etx_passthrough_pending = 0 "Asserted if etx status passthrough is pending - we detected a toggle and have not forwarded the status yet";
    clocked t_sync sync_etx_status_fifo_toggle = {metastable=0, stable=0, last=0};
    comb bit etx_status_fifo_toggle_detected;

    /*b Etx passthrough logic
     */
    etx_passthrough "ETX passthrough logic":
        {
            sync_etx_status_fifo_toggle.metastable <= etx_status_fifo_toggle;
            sync_etx_status_fifo_toggle.stable <= sync_etx_status_fifo_toggle.metastable;
            sync_etx_status_fifo_toggle.last <= sync_etx_status_fifo_toggle.stable;
            etx_status_fifo_toggle_detected = sync_etx_status_fifo_toggle.last ^ sync_etx_status_fifo_toggle.stable;

            if (etx_status_fifo_toggle_detected)
            {
                status_etx_passthrough_pending <= 1;
            }
            if (status_write_passthrough)
            {
                status_etx_passthrough_pending <= 0;
            }
        }

    /*b Registers? Needs new documentation 
     */
    registers "I/O registers and data fifo interface":
        {
            r_mii_rx_data <= mii_data;
            r_mii_rx_dv <= mii_dv;
            r_mii_rx_err <= mii_err;

            next_data_register[4; 0] = data_register[4; 4];
            next_data_register[4; 4] = r_mii_rx_data;
            next_data_register[4; 8] = data_register[4;12];
            next_data_register[4;12] = data_register[4; 0];
            next_data_register[4;16] = data_register[4;20];
            next_data_register[4;20] = data_register[4; 8];
            next_data_register[4;24] = data_register[4;28];
            next_data_register[4;28] = data_register[4;16];

            data_register <= next_data_register;

            if (word_complete)
            {
                data_fifo_data <= next_data_register;
                data_fifo_toggle <= ~data_fifo_toggle;
            }
        }

    /*b Status FIFO interface
     */
    status_fifo_interface "Status FIFO interface":
        {
            status_write_passthrough = 0;
            if ((!status_block_etx_passthrough) && (status_etx_passthrough_pending))
            {
                status_write_passthrough = 1;
            }

            if (status_write || status_write_passthrough)
            {
                status_fifo_toggle <= ~status_fifo_toggle;
                if (status_write_passthrough)
                {
                    status_being_written <= status_to_write_etx_passthrough;
                }
                else
                {
                    status_being_written <= status_to_write;
                }
                status_wait <= 7;
            }
            if (status_wait!=0)
            {
                status_wait <= status_wait-1;
            }
            status_fifo_data = 0;
            status_fifo_data[io_eth_rx_block_byte_length_bits; io_eth_rx_sfd_block_byte_length_start_bit] = 0;
            status_fifo_data[6; io_eth_rx_sfd_block_byte_length_start_bit] = data_fsm.bytes_in_block;
            status_fifo_data[io_eth_rx_packet_byte_length_bits; io_eth_rx_sfd_packet_length_start_bit] = 0;
            status_fifo_data[6; io_eth_rx_sfd_packet_length_start_bit] = data_fsm.bytes_in_block;
            status_fifo_data[10; io_eth_rx_sfd_packet_length_start_bit+6] = data_fsm.blocks_in_packet;
            full_switch (status_being_written)
                {
                case status_to_write_block: // Only mid-packet; always have received 64 bytes!, and the state in data_fsm is unstable and so should be blocked from status FIFO
                {
                    status_fifo_data[io_eth_rx_block_byte_length_bits; io_eth_rx_sfd_block_byte_length_start_bit] = 64;
                    status_fifo_data[6; io_eth_rx_sfd_packet_length_start_bit] = 0;
                    status_fifo_data[io_eth_rx_block_status_bits; io_eth_rx_sfd_block_status_start_bit] = io_eth_rx_status_block_complete;
                }
                case status_to_write_packet_fcs_bad: // At end of packet; guaranteed to have stable bytes_in_block and blocks_in_packet
                {
                    status_fifo_data[io_eth_rx_block_status_bits; io_eth_rx_sfd_block_status_start_bit] = io_eth_rx_status_packet_complete_fcs_bad;
                }
                case status_to_write_packet_fcs_ok: // At end of packet; guaranteed to have stable bytes_in_block and blocks_in_packet
                {
                    status_fifo_data[io_eth_rx_block_status_bits; io_eth_rx_sfd_block_status_start_bit] = io_eth_rx_status_packet_complete_fcs_ok;
                }
                case status_to_write_fifo_overrun: // At end of packet; guaranteed to have stable bytes_in_block and blocks_in_packet
                {
                    status_fifo_data[io_eth_rx_block_status_bits; io_eth_rx_sfd_block_status_start_bit] = io_eth_rx_status_fifo_overrun;
                }
                case status_to_write_odd_nybbles: // At end of packet; guaranteed to have stable bytes_in_block and blocks_in_packet
                {
                    status_fifo_data[io_eth_rx_block_status_bits; io_eth_rx_sfd_block_status_start_bit] = io_eth_rx_status_packet_complete_odd_nybbles;
                }
                case status_to_write_rx_err:
                {
                    status_fifo_data[io_eth_rx_block_status_bits; io_eth_rx_sfd_block_status_start_bit] = io_eth_rx_status_block_complete;
                }
                case status_to_write_etx_passthrough:
                {
                    status_fifo_data = etx_status_fifo_data;
                    status_fifo_data[31] = 1;
                }
                }
    }

    /*b Data FSM, block_complete and word_complete indications; block_complete is a subset of word_complete
     */
    data_fsm "Data FSM":
        {
            next_data_fsm = {state=data_fsm.state, bytes_in_block=data_fsm.bytes_in_block, counter=data_fsm.counter+1, blocks_in_packet=data_fsm.blocks_in_packet};
            data_fsm <= next_data_fsm;
            word_complete = 0;
            status_write <= 0;
            status_block_etx_passthrough = (status_wait!=0);
            full_switch (data_fsm.state)
                {
                case data_fsm_idle: // if there is good data then start receiving it; if there is bad data then its a framing error; do not block etx status pass-through
                {
                    next_data_fsm.counter = 0;
                    if ( r_mii_rx_dv )
                    {
                        if (r_mii_rx_err)
                        {
                            next_data_fsm.state = data_fsm_framing_error;
                        }
                        elsif (r_mii_rx_data==4h5) // Preamble
                            {
                                next_data_fsm.state = data_fsm_wait_for_end_of_sfd;
                            }
                        else
                        {
                            next_data_fsm.state = data_fsm_idle;
                        }
                    }
                }
                case data_fsm_wait_for_end_of_sfd: // if there is more sfd then stay, else end of sfd then start receiving data with appropriate padding skip; do not block etx status pass-through
                {
                    next_data_fsm.counter = 0;
                    next_data_fsm.bytes_in_block = 0;
                    next_data_fsm.blocks_in_packet = 0;
                    full_switch (cfg_padding)
                    {
                    case 0:
                    {
                        next_data_fsm.counter = 0;
                        next_data_fsm.bytes_in_block = 0;
                    }
                    case 1:
                    {
                        next_data_fsm.counter = 2;
                        next_data_fsm.bytes_in_block = 1;
                    }
                    case 2:
                    {
                        next_data_fsm.counter = 4;
                        next_data_fsm.bytes_in_block = 2;
                    }
                    case 3:
                    {
                        next_data_fsm.counter = 6;
                        next_data_fsm.bytes_in_block = 3;
                    }
                    }
                    if ( r_mii_rx_dv )
                    {
                        if (r_mii_rx_err)
                        {
                            next_data_fsm.state = data_fsm_framing_error;
                        }
                        elsif (r_mii_rx_data==4h5) // Preamble
                            {
                                next_data_fsm.state = data_fsm_wait_for_end_of_sfd;
                            }
                        elsif (r_mii_rx_data==4hd) // SFD
                            {
                                next_data_fsm.state = data_fsm_reading_data;
                            }
                        else
                        {
                            next_data_fsm.state = data_fsm_idle;
                        }
                    }
                    else
                    {
                        next_data_fsm.state = data_fsm_idle;
                    }
                }
                case data_fsm_reading_data: // read data until last nybble received, but handle next-to-last nybble of word by punting; block etx status pass-through if we are near the end of a block
                {
                    if (data_fsm.bytes_in_block[3;3]==7) // if there are 56 to 63 bytes in our current block then block the etx passthrough
                    {
                        status_block_etx_passthrough = 1;
                    }
                    if ( !r_mii_rx_dv )
                    {
                        if (data_fsm.counter[0]==0)
                        {
                            next_data_fsm.state = data_fsm_packet_complete_waiting; // Don't reset count - we want to wait in the next state until counter[4;0]==0 (i.e. 1 to 7 cycles)
                            status_to_write <= fcs_ok ? status_to_write_packet_fcs_bad : status_to_write_packet_fcs_ok;
                        }
                        else // Data valid taken away mid-byte
                        {
                            next_data_fsm.counter = 0;
                            next_data_fsm.state = data_fsm_framing_error;
                            status_to_write <= status_to_write_odd_nybbles;
                        }
                    }
                    else
                    {
                        if ( r_mii_rx_err ) // Error in the nybble
                        {
                            next_data_fsm.counter = 0;
                            next_data_fsm.state = data_fsm_framing_error;
                            status_to_write <= status_to_write_rx_err;
                        }
                        else
                        {
                            if (data_fsm.counter[0]==1)
                            {
                                next_data_fsm.bytes_in_block = data_fsm.bytes_in_block+1;
                            }
                            if (data_fsm.counter==6) // Last nybble of a word coming next
                            {
                                next_data_fsm.state = data_fsm_reading_data_last_nybble_of_word;
                            }
                        }
                    }
                }
                case data_fsm_reading_data_last_nybble_of_word: // 7th nybble of a word should be ready; if not we have a framing error, if we do write the word and a status if we hit the 16th word
                {
                    if (data_fsm.bytes_in_block[3;3]==7) // if there are 56 to 63 bytes in our current block then block the etx passthrough
                    {
                        status_block_etx_passthrough = 1;
                    }
                    next_data_fsm.counter = 0;
                    if ( !r_mii_rx_dv ) // Data valid taken away mid-byte
                    {
                        next_data_fsm.state = data_fsm_framing_error;
                        status_to_write <= status_to_write_odd_nybbles;
                    }
                    else
                    {
                        if ( r_mii_rx_err ) // Error in the nybble
                        {
                            next_data_fsm.state = data_fsm_framing_error;
                            status_to_write <= status_to_write_rx_err;
                        }
                        elsif (data_fifo_full)
                            {
                                assert(0,"Ethernet receive data fifo full");
                                next_data_fsm.counter = 0;
                                next_data_fsm.state = data_fsm_framing_error;
                                status_to_write <= status_to_write_fifo_overrun;
                            }
                        else
                        {
                            next_data_fsm.bytes_in_block = data_fsm.bytes_in_block+1;
                            next_data_fsm.state = data_fsm_reading_data;
                            word_complete = 1;
                            if (next_data_fsm.bytes_in_block==0) // Read a whole block - tell the status FIFO
                            {
                                next_data_fsm.blocks_in_packet = data_fsm.blocks_in_packet+1;
                                status_to_write <= status_to_write_block;
                                status_write <= 1;
                            }
                        }
                    }
                }
                case data_fsm_packet_complete_waiting: // Shifting the data up - guarantees a gap between last word write/block write and next one, also; we sit in here for from 1 to 7 cycles
                {
                    // there will be enough time before the complete status goes, so we do not need to block etx status passthrough
                    if (data_fsm.counter == 7)
                    {
                        next_data_fsm.state = data_fsm_packet_complete;
                        if (data_fsm.bytes_in_block[2;0]!=0)
                        {
                            word_complete = 1; // Data will have been shifted up to top nybble during the waiting state; but there is no word if we were given a precise word-length packet. Hm.
                        }
                    }
                }
                case data_fsm_packet_complete: // Always entered with counter of 0. Wrote a whole packet except last word; write last word (if any bytes ready) and write status giving full status of packet
                {
                    status_block_etx_passthrough = 1; // there will not be enough time
                    if (data_fsm.counter==7)
                    {
                        next_data_fsm.state = data_fsm_idle;
                        status_write <= 1; // Guaranteed to be 8 cycles or more from last block_complete or etx passthrough
                    }
                }
                case data_fsm_framing_error: // Framing error; we enter with counter of 0, and wait for 8 cycles, then we present a status. Wait for status and data FIFO to complete any pending writes, then write last word (if any bytes ready) and write status
                {
                    if (r_mii_rx_dv)
                    {
                        next_data_fsm.counter = 0;
                        // there will be enough time from here to our framing error status write since we reset the counter here - so dont block etx passthrough
                    }
                    else
                    {
                        status_block_etx_passthrough = 1; // there will not be enough time if dv stays away, so block passthrough
                        if (data_fsm.counter == 7)
                        {
                            next_data_fsm.state = data_fsm_idle;
                            status_write <= 1; // Guaranteed to be 8 cycles or more from last block_complete, and we will be in idle before (at worst) hitting framing error again, eight cycles prior to status write
                        }
                    }
                }
                }
        }

    /*b FCS calculation - fcs, next_fcs, data_for_fcs, fcs_ok
     */
    fcs "Calculate FCS from transmit nybbles":
        {
            next_fcs[4;0] = 0;
            next_fcs[28;4] = fcs[28;0];
            data_for_fcs[0] = fcs[31] ^ r_mii_rx_data[0]; // Bit 0 is the first on the wire, so it goes with bit 31 of the FCS
            data_for_fcs[1] = fcs[30] ^ r_mii_rx_data[1]; // Bit 1 comes next, so it takes bit 30 of FCS
            data_for_fcs[2] = fcs[29] ^ r_mii_rx_data[2]; // etc
            data_for_fcs[3] = fcs[28] ^ r_mii_rx_data[3];
            if (data_for_fcs[3])
            {
                next_fcs = next_fcs ^ 32b00000100110000010001110110110111; // poly is 32.26.23.22.16.12.11.10.8.7.5.4.2.1.0
            }
            if (data_for_fcs[2])
            {
                next_fcs = next_fcs ^ 32b00001001100000100011101101101110; // rotate in one bit
            }
            if (data_for_fcs[1])
            {
                next_fcs = next_fcs ^ 32b00010011000001000111011011011100; // rotate in two bits
            }
            if (data_for_fcs[0])
            {
                next_fcs = next_fcs ^ 32b00100110000010001110110110111000; // rotate in three bits
            }

            fcs <= 32hffffffff;
            part_switch (data_fsm.state)
                {
                case data_fsm_reading_data:
                {
                    fcs <= next_fcs;
                }
                case data_fsm_packet_complete_waiting:
                {
                    fcs <= fcs;
                }
                }
            fcs_ok = (fcs==32hc704dd7b);
        }

    /*b All done
     */
}
