/*a Includes
 */
include "postbus.h"

/*a Types
 */
/*t t_arb_fsm
 */
typedef fsm
{
    arb_fsm_idle;
    arb_fsm_src_0;
    arb_fsm_src_1;
    arb_fsm_src_2;
    arb_fsm_src_3;
} t_arb_fsm;

/*a postbus_input_mux module
 */
module postbus_input_mux( input clock int_clock, input bit int_reset,
                          input t_postbus_type src_type_0, input t_postbus_data src_data_0, output t_postbus_ack src_ack_0,
                          input t_postbus_type src_type_1, input t_postbus_data src_data_1, output t_postbus_ack src_ack_1,
                          input t_postbus_type src_type_2, input t_postbus_data src_data_2, output t_postbus_ack src_ack_2,
                          input t_postbus_type src_type_3, input t_postbus_data src_data_3, output t_postbus_ack src_ack_3,
                          input t_postbus_ack tgt_ack, output t_postbus_type tgt_type,
                          output t_postbus_data tgt_data
    )
    "This is a 4-to-1 postbus multiplexer, which is designed as the input source to a
    registering 1-to-n postbus multiplexer";
{
    /*b State and combinatorials
     */
    clocked rising int_clock active_high int_reset t_arb_fsm state = arb_fsm_idle;
    clocked rising int_clock active_high int_reset bit src_first_word = 0 "High if the source is presenting the first word of a transaction";
    comb t_arb_fsm next_state "Next state of FSM";
    comb bit wait "Set if a transfer is in place and the selected target indicates no acknowledge";

    /*b Arbitration FSM - state, next_state, wait
     */
    fsm "Arbitration FSM  - select next source to transfer; this is more complex than it need be, as it allows for back-to-back transfers from different masters.":
        {
            next_state = state;
            wait = 0;
            if (state!=arb_fsm_idle)
            {
                wait = tgt_ack;
            }
            full_switch (state)
                {
                case arb_fsm_idle:
                    if (src_type_3==postbus_word_type_start) { next_state = arb_fsm_src_3; }
                    if (src_type_2==postbus_word_type_start) { next_state = arb_fsm_src_2; }
                    if (src_type_1==postbus_word_type_start) { next_state = arb_fsm_src_1; }
                    if (src_type_0==postbus_word_type_start) { next_state = arb_fsm_src_0; }
                case arb_fsm_src_0:
                    if ( (src_type_0==postbus_word_type_last) || ((src_first_word) && (src_data_0[0])) )
                    {
                        next_state = arb_fsm_idle;
                        if (src_type_3==postbus_word_type_start) { next_state = arb_fsm_src_3; }
                        if (src_type_2==postbus_word_type_start) { next_state = arb_fsm_src_2; }
                        if (src_type_1==postbus_word_type_start) { next_state = arb_fsm_src_1; }
                    }
                case arb_fsm_src_1:
                    if ( (src_type_1==postbus_word_type_last) || ((src_first_word) && (src_data_1[0])) )
                    {
                        next_state = arb_fsm_idle;
                        if (src_type_0==postbus_word_type_start) { next_state = arb_fsm_src_0; }
                        if (src_type_3==postbus_word_type_start) { next_state = arb_fsm_src_3; }
                        if (src_type_2==postbus_word_type_start) { next_state = arb_fsm_src_2; }
                    }
                case arb_fsm_src_2:
                    if ( (src_type_2==postbus_word_type_last) || ((src_first_word) && (src_data_2[0])) )
                    {
                        next_state = arb_fsm_idle;
                        if (src_type_1==postbus_word_type_start) { next_state = arb_fsm_src_1; }
                        if (src_type_0==postbus_word_type_start) { next_state = arb_fsm_src_0; }
                        if (src_type_3==postbus_word_type_start) { next_state = arb_fsm_src_3; }
                    }
                case arb_fsm_src_3:
                    if ( (src_type_3==postbus_word_type_last) || ((src_first_word) && (src_data_3[0])) )
                    {
                        next_state = arb_fsm_idle;
                        if (src_type_2==postbus_word_type_start) { next_state = arb_fsm_src_2; }
                        if (src_type_1==postbus_word_type_start) { next_state = arb_fsm_src_1; }
                        if (src_type_0==postbus_word_type_start) { next_state = arb_fsm_src_0; }
                    }
                }
            if (wait)
            {
                next_state = state;
            }
            state <= next_state;
        }

    /*b Determine first cycle of a transaction - src_first_word
     */
    first_of_transaction "Determine first cycle of a transaction":
        {
            if (next_state != state)
            {
                src_first_word <= 1;
            }
            else
            {
                if (!wait)
                {
                    src_first_word <= 0;
                }
            }
        }

    /*b Output muxes for data and target - tgt_data, tgt_type
     */
    output_mux "Output data, type multiplexers":
        {
            full_switch(state)
                {
                case arb_fsm_idle:
                    tgt_data = src_data_0;
                    tgt_type = postbus_word_type_idle;
                case arb_fsm_src_0: 
                    tgt_data = src_data_0;
                    tgt_type = src_type_0;
                case arb_fsm_src_1: 
                    tgt_data = src_data_1;
                    tgt_type = src_type_0;
                case arb_fsm_src_2: 
                    tgt_data = src_data_2;
                    tgt_type = src_type_0;
                case arb_fsm_src_3: 
                    tgt_data = src_data_3;
                    tgt_type = src_type_0;
                }
        }

    /*b Drive selected acknowledge - src_ack_*
     */
    ack_drive "Acknowledge drivers":
        {
            src_ack_0 = 0;
            src_ack_1 = 0;
            src_ack_2 = 0;
            src_ack_3 = 0;
            part_switch(state)
                {
                case arb_fsm_src_0: src_ack_0 = tgt_ack;
                case arb_fsm_src_1: src_ack_1 = tgt_ack;
                case arb_fsm_src_2: src_ack_2 = tgt_ack;
                case arb_fsm_src_3: src_ack_3 = tgt_ack;
                }
        }
}
