/*a Includes
 */
include "gip.h"
include "gip_internal.h"

/*a External modules
 */
/*m gip_alu_arith_op_data_path
 */
extern module gip_alu_arith_op_data_path( input t_gip_word op_a,
                                   input bit zero_a,
                                   input bit negate_a,
                                   input t_gip_word op_b,
                                   input bit zero_b,
                                   input bit negate_b,
                                   input bit use_shifted_b,
                                   input bit c_in,
                                   output t_gip_word sum,
                                   output bit z_out,
                                   output bit n_out,
                                   output bit c_out,
                                   output bit v_out )
{
    timing comb input op_a, zero_a, negate_a;
    timing comb input op_b, zero_b, negate_b, use_shifted_b;
    timing comb input c_in;
    timing comb output sum;
    timing comb output z_out, n_out, c_out, v_out;
}


/*a Modules
 */
module gip_alu_arith_op( input t_gip_word op_a,
                         input t_gip_word op_b,
                         input bit c_in,
                         input bit p_in,
                         input bit[2] shf,
                         input t_gip_arith_op arith_op,
                         output t_gip_word result,
                         output bit z,
                         output bit n,
                         output bit v,
                         output bit c,
                         output bit shf_carry_override,
                         output bit shf_carry_out )
"
This module implements the arithmetic operations for the GIP
"
{
    comb bit zero_a;
    comb bit negate_a;
    comb bit zero_b;
    comb bit negate_b;
    comb bit use_shifted_b;
    comb bit dp_c_in;
    net t_gip_word sum;
    net bit dp_z_out;
    net bit dp_n_out;
    net bit dp_c_out;
    net bit dp_v_out;
   
    /*b Determine adder inputs
     */
    adder_inputs "Determine adder inputs from instruction and multiply state":
        {
            shf_carry_override = 0;
            shf_carry_out = 0;
            dp_c_in = 0;
            zero_a = 0;
            negate_a = 0;
            zero_b = 0;
            negate_b = 0;
            use_shifted_b = 0;

            part_switch (arith_op)
            {
            case gip_arith_op_add:
            {
                dp_c_in = 0;
            }
            case gip_arith_op_adc:
            {
                dp_c_in = c_in;
            }
            case gip_arith_op_sub:
            {
                negate_b = 1;
                dp_c_in = 1;
            }
            case gip_arith_op_sbc:
            {
                negate_b = 1;
                dp_c_in = 1;
            }
            case gip_arith_op_rsub:
            {
                negate_a = 1;
                dp_c_in = 1;
            }
            case gip_arith_op_rsbc:
            {
                negate_a = 1;
                dp_c_in = c_in;
            }
            case gip_arith_op_init:
            {
                zero_a = 1;
                dp_c_in = 0;
            }
            case gip_arith_op_mla:
            case gip_arith_op_mlb:
            {
                zero_b = 1;
                shf_carry_override = 1;
                if (p_in)
                {
                    full_switch (shf)
                    {
                    case 0:{ zero_b = 0;        dp_c_in=0; shf_carry_out=0; } // net mult by 1   => +b
                    case 1:{ use_shifted_b = 1; dp_c_in=0; shf_carry_out=0; } // net mult by 2   => +2b
                    case 2:{ negate_b = 1;      dp_c_in=1; shf_carry_out=1; } // net mult by 4-1 => +3b
                    case 3:{ zero_b=1;          dp_c_in=0; shf_carry_out=1; } // net mult by 4   => +4b
                    }
                }
                else
                {
                    full_switch (shf)
                    {
                    case 0:{ zero_b = 1;        dp_c_in=0; shf_carry_out=0; } // net mult by 0   => +0
                    case 1:{ zero_b = 0;        dp_c_in=0; shf_carry_out=0; } // net mult by 1   => +b
                    case 2:{ use_shifted_b = 1; dp_c_in=0; shf_carry_out=0; } // net mult by 2   => +2b
                    case 3:{ negate_b = 1;      dp_c_in=1; shf_carry_out=1; } // net mult by 4-1 => +3b
                    }
                }
            }
            }
        }

    /*b Adder datapath
     */
    adder_datapath "Adder datapath":
        {
            gip_alu_arith_op_data_path data_path( op_a <= op_a,
                                                  op_b <= op_b,
                                                  zero_a <= zero_a,
                                                  negate_a <= negate_a,
                                                  zero_b <= zero_b,
                                                  negate_b <= negate_b,
                                                  use_shifted_b <= use_shifted_b,
                                                  c_in <= dp_c_in,
                                                  sum => sum,
                                                  z_out => dp_z_out,
                                                  n_out => dp_n_out,
                                                  c_out => dp_c_out,
                                                  v_out => dp_v_out );

        }

    /*b Final result
     */
    final_result "Final result selection/operation":
        {
            z = dp_z_out;
            n = dp_n_out;
            c = dp_c_out;
            v = dp_v_out;
            if (arith_op==gip_arith_op_write_flags)
            {
                z = op_b[0];
                n = op_b[1];
                c = op_b[2];
                v = op_b[3];
            }
            result = sum;
        }

    /*b Done
     */
}
