/*a Copyright Gavin J Stark, 2004
 */

/*a Includes
 */
include "io_uart.h"

/*a Types
 */

/*a External modules required
 */
/*m apb_target_uart
 */
extern module apb_target_ext_bus_master( clock apb_clock "Internal system clock",
                                  input bit int_reset "Internal reset",

                                  input bit[3] apb_paddr,
                                  input bit apb_penable,
                                  input bit apb_pselect,
                                  input bit[32] apb_pwdata,
                                  input bit apb_prnw,
                                  output bit[32] apb_prdata,
                                  output bit apb_pwait,

                                  output bit[4]ext_bus_ce,
                                  output bit ext_bus_oe,
                                  output bit ext_bus_we,
                                  output bit[24]ext_bus_address,
                                  output bit ext_bus_write_data_enable,
                                  output bit[32]ext_bus_write_data,
                                  input bit[32]ext_bus_read_data
                                  )
{
    timing to rising clock apb_clock int_reset;

    timing to rising clock apb_clock apb_pselect, apb_penable, apb_paddr, apb_pwdata, apb_prnw;
    timing comb input apb_pselect, apb_penable, apb_paddr, apb_prnw;
    timing from rising clock apb_clock apb_prdata;
    timing comb output apb_prdata;

    timing to rising clock apb_clock ext_bus_read_data;
    timing from rising clock apb_clock ext_bus_ce, ext_bus_oe, ext_bus_we, ext_bus_address, ext_bus_write_data_enable, ext_bus_write_data;
}

/*m apb_target_uart
 */
extern module apb_target_uart( clock apb_clock "Internal system clock",
                         input bit int_reset "Internal reset",

                         input bit[3] apb_paddr,
                         input bit apb_penable,
                         input bit apb_pselect,
                         input bit[32] apb_pwdata,
                         input bit apb_prnw,
                        output bit[32] apb_prdata,

                         output bit cmd_fifo_empty,
                         output bit[32] cmd_fifo_data,
                         input bit cmd_fifo_toggle,

                         output bit status_fifo_full,
                         input bit status_fifo_toggle,
                         input bit[32] status_fifo_data )
{
    timing to rising clock apb_clock int_reset;

    timing to rising clock apb_clock apb_pselect, apb_penable, apb_paddr, apb_pwdata, apb_prnw;
    timing comb input apb_pselect, apb_penable, apb_paddr, apb_prnw;
    timing from rising clock apb_clock apb_prdata;
    timing comb output apb_prdata;

    timing to rising clock apb_clock cmd_fifo_toggle;
    timing from rising clock apb_clock cmd_fifo_empty, cmd_fifo_data;
    timing to rising clock apb_clock status_fifo_toggle, status_fifo_data;
    timing from rising clock apb_clock status_fifo_full;
}

/*a Modules
 */
module apb_devices( clock int_clock,
                    input bit int_reset,

                    input bit apb_pselect,
                    input bit apb_penable,
                    input bit apb_prnw,
                    input bit[5] apb_paddr,
                    input bit[32] apb_pwdata,
                    output bit[32] apb_prdata,
                    output bit apb_pwait,

                    input bit[8] switches,
                    output bit[8] leds,
                    output bit txd,
                    input bit rxd,
                    output bit[4]ext_bus_ce,
                    output bit ext_bus_oe,
                    output bit ext_bus_we,
                    output bit[24]ext_bus_address,
                    output bit ext_bus_write_data_enable,
                    output bit[32]ext_bus_write_data,
                    input bit[32]ext_bus_read_data
    )
{
    default clock int_clock;
    default reset int_reset;

//    comb bit[8] leds;
    net bit txd;

    net bit[4]ext_bus_ce;
    net bit ext_bus_oe;
    net bit ext_bus_we;
    net bit[24]ext_bus_address;
    net bit ext_bus_write_data_enable;
    net bit[32]ext_bus_write_data;

    clocked bit[24] clock_divider=0;
    comb bit clock_enable;

    comb bit tx_baud_enable "Baud enable for transmit, 16 x bit time";
//    net bit txd "Transmit data out";
//    net bit txd_fc "Transmit flow control; assert to pause transmit";

    comb bit rx_baud_enable "Baud enable for receive, 16 x bit time";
//    net bit rxd "Receive data in";
    net bit rxd_fc "Receive flow control; asserted to pause transmit";

    net bit cmd_fifo_empty;
    net bit[32] cmd_fifo_data;
    net bit cmd_fifo_toggle;

    net bit status_fifo_full;
    net bit status_fifo_toggle;
    net bit[32] status_fifo_data;

//    net bit[32] apb_prdata;
    net bit[32] apb_prdata_uart;
    net bit[32] apb_prdata_ext_bus;
    net bit apb_pwait;

    comb bit[2] cfg_uart_speed;
    comb bit[16] cfg_baud_divider;
    clocked bit[16] baud_counter=0;
    clocked bit toggle=0;
    clocked bit[6] baud_divider = 0;
    clocked bit toggle_2=0;

    /*b Clock divider
     */
    divider "Clock divider for LED":
        {
            cfg_uart_speed = switches[2;0];
            clock_divider <= clock_divider+1;
            clock_enable = 0;
            if ((clock_divider[8;12]==switches) && (clock_divider[12;0]==0))
//            if (clock_divider[10;0]==0)
            {
                toggle <= ~toggle;
                clock_enable = 1;
                clock_divider <= 0;
            }
            leds = clock_divider[8;11];
            leds[0] = toggle;
            leds[1] = toggle_2;
            leds[2] = txd;
            leds[3] = rxd;
            full_switch( cfg_uart_speed )
                {
                case 0: // 260=>9600 - actually 1200 for 5MHz; for 125/12 we need 60
                {
                    cfg_baud_divider = 260;
                    cfg_baud_divider = 68;
                }
                case 1: // 130=>19200 - actually 2400 for 5MHz and for 125/12 we need 241
                {
                    cfg_baud_divider = 130;
                    cfg_baud_divider = 271;
                }
                case 2: // 38400 - NOW 10Hz for 5MHz
                {
                    cfg_baud_divider = 65;
                    cfg_baud_divider = 16h7a21; // 31250 = 5,000,000/160
                    cfg_baud_divider = 34;
                }
                case 3: // none - i.e. divide by 8
                {
                    cfg_baud_divider = 8;
                }
                }
            baud_counter <= baud_counter+1;
            if (baud_counter+1 == cfg_baud_divider)
            {
                baud_counter <= 0;
            }
            rx_baud_enable = (baud_counter==0);
            tx_baud_enable = rx_baud_enable;
            if (rx_baud_enable)
            {
                baud_divider <= baud_divider+1;
                if (baud_divider==0)
                {
                    toggle_2 <= ~toggle_2;
                }
            }
        }

    /*b APB instances
     */
    apb_instances "APB Instances":
        {
            apb_target_ext_bus_master ext_bus_apb( apb_clock <- int_clock,
                                                   int_reset <= int_reset,

                                                   apb_pselect <= apb_pselect && (apb_paddr[2;3]==1),
                                                   apb_penable <= apb_penable,
                                                   apb_paddr <= apb_paddr[3;0],
                                                   apb_prnw <= apb_prnw,
                                                   apb_pwdata <= apb_pwdata,
                                                   apb_prdata => apb_prdata_ext_bus,
                                                   apb_pwait => apb_pwait,

                                                   ext_bus_ce => ext_bus_ce,
                                                   ext_bus_oe => ext_bus_oe,
                                                   ext_bus_we => ext_bus_we,
                                                   ext_bus_address => ext_bus_address,
                                                   ext_bus_write_data_enable => ext_bus_write_data_enable,
                                                   ext_bus_write_data => ext_bus_write_data,
                                                   ext_bus_read_data <= ext_bus_read_data );


            apb_target_uart uart_apb( apb_clock <- int_clock,
                                      int_reset <= int_reset,

                                      apb_pselect <= apb_pselect && (apb_paddr[2;3]==0),
                                      apb_penable <= apb_penable,
                                      apb_paddr <= apb_paddr[3;0],
                                      apb_prnw <= apb_prnw,
                                      apb_pwdata <= apb_pwdata,
                                      apb_prdata => apb_prdata_uart,
                                      
                                      cmd_fifo_empty => cmd_fifo_empty,
                                      cmd_fifo_data => cmd_fifo_data,
                                      cmd_fifo_toggle <= cmd_fifo_toggle,

                                      status_fifo_full => status_fifo_full,
                                      status_fifo_data <= status_fifo_data,
                                      status_fifo_toggle <= status_fifo_toggle );

            io_uart uart_io( int_clock <- int_clock,
                          int_reset <= int_reset,
                          tx_baud_enable <= tx_baud_enable,
                          txd => txd,
                          txd_fc <= 0,
                          rx_baud_enable <= rx_baud_enable,
                          rxd <= rxd | switches[2],
                          rxd_fc => rxd_fc,

                          cmd_fifo_empty <= cmd_fifo_empty,
                          cmd_fifo_data <= cmd_fifo_data,
                          cmd_fifo_toggle => cmd_fifo_toggle,

                          status_fifo_full <= status_fifo_full,
                          status_fifo_data => status_fifo_data,
                          status_fifo_toggle => status_fifo_toggle );

            apb_prdata = (apb_paddr[2;3]==0)?apb_prdata_uart : apb_prdata_ext_bus;
        }

}

