/*a Copyright Gavin J Stark, 2004
 */

/*a To do
 */

/*a Constants
 */

/*a Types
 */
/*t t_sync_toggle
 */
typedef struct {
    bit[2] sync;
    bit last;
} t_sync_toggle;

/*a fifo_ctrl_synch
 */
module fifo_ctrl_synch( clock int_clock,
                        input bit int_reset,
                        input bit valid_in "Valid signal from the I/O clock domain; synchronized and edge detected for a request",
                        output bit request "Internal clock domain signal, asserted and deasserted synchronously",
                        input bit acknowledge "Internal clock domain signal, combinatorially generated from requests; indicates request should be removed in next cycle" )

    /*b Documentation
     */
    "
This module implements the simple synchronized command and request validation scheme used with the I/O FIFOs.

A single signal from the I/O clock domain is synchronized and edge-detected.

An edge indicates that the request the I/O system is presenting is valid; this subsystem detects that and presents the request, which is removed when the request is acknowledged.

There is no handshake back to the I/O clock domain; the internal clock domain is responsible for handling the requests presented within strict guarantees for each I/O device, making the handshake unnecessary.

"
{

    /*b Clock and reset
     */
    default clock int_clock;
    default reset int_reset;

    /*b Synchronizer
     */
    clocked t_sync_toggle sync_toggle = { sync=0, last = 0 } "Synchronizer";
    comb bit toggled "Indication that the synchronizer has toggled";
    clocked bit request_pending=0 "Asserted if a request is pending; that is if it has been presented once, but has not been acknowledged";

    /*b Synchronizer code
     */
    synchronizer "Synchronizer code":
        {
            sync_toggle.sync[0] <= valid_in;
            sync_toggle.sync[1] <= sync_toggle.sync[0];
            sync_toggle.last    <= sync_toggle.sync[1];

            toggled = (sync_toggle.last!=sync_toggle.sync[1]);
            request = request_pending || toggled;
            if (acknowledge)
            {
                request_pending <= 0;
            }
            else
            {
                request_pending <= request;
            }
        }
}
