/*a Copyright Gavin J Stark, 2004
 */

/*a To do
 */

/*a Includes
 */
include "io_simple_fifo.h"

/*a Types
 */
typedef struct
{
    bit[io_simple_fifo_address_size] read_ptr;
    bit[io_simple_fifo_address_size] write_ptr;

    bit empty;
    bit full;
    bit watermark;
    bit overflowed;
    bit underflowed;
} t_fifo_state;

typedef struct
{
    bit[io_simple_fifo_address_size] base_address;
    bit[io_simple_fifo_address_size] size_m_one;
    bit[io_simple_fifo_address_size] watermark;
} t_fifo_cfg;

/*a Module
 */
module io_simple_fifo( clock int_clock "main system clck",
                              input bit int_reset "main system reset",
                              input t_simple_fifo_op fifo_op "Operation to perform",
                              output bit[io_simple_fifo_address_size] fifo_write_address "Write address out",
                              output bit[io_simple_fifo_address_size] fifo_read_address "Read address out",

                              output bit fifo_empty "Asserted if more than zero entries are present",
                              output bit fifo_watermark "Asserted if more than 'watermark' entries are present",
                              output bit fifo_full "Asserted if read_ptr==write_ptr and not empty",
                              output bit fifo_overflowed "Asserted if the FIFO has overflowed since last reset or configuration write",
                              output bit fifo_underflowed  "Asserted if the FIFO has underflowed since last reset or configuration write",

                              input bit[io_simple_fifo_address_size] cfg_base_address,
                              input bit[io_simple_fifo_address_size] cfg_size_m_one,
                              input bit[io_simple_fifo_address_size] cfg_watermark )
{
    default clock int_clock;
    default reset int_reset;

    comb bit inc_read_ptr;
    comb bit inc_write_ptr;
    comb t_fifo_state next_fifo_state;
    comb bit[io_simple_fifo_address_size] current_entries;
    comb bit[io_simple_fifo_address_size] next_entries;

    clocked t_fifo_state fifo_state = { empty=1,
                                        full=0, 
                                        watermark=0,
                                        overflowed=0,
                                        underflowed=0,
                                        read_ptr=0,
                                        write_ptr=0 };
    clocked t_fifo_cfg fifo_cfg = { base_address=0, size_m_one=0, watermark=0 };

    fifo_outputs "Drive the outputs":
        {
            fifo_write_address = fifo_cfg.base_address + fifo_state.write_ptr;
            fifo_read_address  = fifo_cfg.base_address + fifo_state.read_ptr;

            fifo_empty = fifo_state.empty;
            fifo_full = fifo_state.full;
            fifo_watermark = fifo_state.watermark;
            fifo_overflowed = fifo_state.overflowed;
            fifo_underflowed = fifo_state.underflowed;
        }

    next_fifo "Determine next state of FIFO if incrementing either ptr":
        {
            
            next_fifo_state = fifo_state;
            next_entries = current_entries;
            if (inc_write_ptr)
            {
                if (fifo_state.full)
                {
                    next_fifo_state.overflowed = 1;
                }
                else
                {
                    if (fifo_state.write_ptr == fifo_cfg.size_m_one)
                    {
                        next_fifo_state.write_ptr = 0;
                    }
                    else
                    {
                        next_fifo_state.write_ptr = fifo_state.write_ptr+1;
                    }
                    next_entries = current_entries+1;
                    next_fifo_state.full = (current_entries==fifo_cfg.size_m_one);
                }
            }
            if (inc_read_ptr)
            {
                if (fifo_state.empty)
                {
                    next_fifo_state.underflowed = 1;
                }
                else
                {
                    if (fifo_state.read_ptr == fifo_cfg.size_m_one)
                    {
                        next_fifo_state.read_ptr = 0;
                    }
                    else
                    {
                        next_fifo_state.read_ptr = fifo_state.read_ptr+1;
                    }
                    next_entries = current_entries-1;
                    next_fifo_state.empty = (next_entries==0);
                }
            }
            next_fifo_state.watermark = next_fifo_state.full | (next_entries>fifo_cfg.size_m_one);
        }

    count_entries "Count number of entries in FIFO":
        {
            current_entries = fifo_state.write_ptr - fifo_state.read_ptr;
            if (fifo_state.write_ptr<fifo_state.read_ptr)
            {
                current_entries = current_entries+fifo_cfg.size_m_one+1;
            }
            if ((fifo_state.write_ptr==fifo_state.read_ptr) && (fifo_state.full))
            {
                current_entries = current_entries+fifo_cfg.size_m_one+1;
            }
        }

    fifo_operation "Handle the FIFO":
        {
            full_switch (fifo_op)
                {
                case simple_fifo_op_write_cfg:
                {
                    fifo_state <= { empty=1, full=0, watermark=0, overflowed=0, underflowed=0, read_ptr=0, write_ptr=0 };
                    fifo_cfg <= { base_address=cfg_base_address, size_m_one=cfg_size_m_one, watermark=cfg_watermark };
                }
                case simple_fifo_op_reset:
                {
                    fifo_state <= { empty=1, full=0, watermark=0, overflowed=0, underflowed=0, read_ptr=0, write_ptr=0 };
                }
                case simple_fifo_op_inc_write_ptr:
                {
                    inc_write_ptr = 1;
                    fifo_state <= next_fifo_state;
                }
                case simple_fifo_op_inc_read_ptr:
                {
                    inc_read_ptr = 1;
                    fifo_state <= next_fifo_state;
                }
                }
        }
}

