include "postbus.h"

typedef fsm
{
    arb_fsm_idle;
    arb_fsm_xfr_0;
    arb_fsm_xfr_1;
    arb_fsm_xfr_2;
    arb_fsm_xfr_3;
} t_arb_fsm;

module simple_postbus_router( clock int_clock, input bit int_reset,
                              input t_postbus_type src_type_0, input t_postbus_data src_data_0, output t_postbus_ack src_ack_0,
                              input t_postbus_type src_type_1, input t_postbus_data src_data_1, output t_postbus_ack src_ack_1,
                              input t_postbus_type src_type_2, input t_postbus_data src_data_2, output t_postbus_ack src_ack_2,
                              input t_postbus_type src_type_3, input t_postbus_data src_data_3, output t_postbus_ack src_ack_3,
                              input t_postbus_ack tgt_ack_0, output t_postbus_type tgt_type_0,
                              input t_postbus_ack tgt_ack_1, output t_postbus_type tgt_type_1,
                              input t_postbus_ack tgt_ack_2, output t_postbus_type tgt_type_2,
                              input t_postbus_ack tgt_ack_3, output t_postbus_type tgt_type_3,
                              input t_postbus_ack tgt_ack_4, output t_postbus_type tgt_type_4,
                              input t_postbus_ack tgt_ack_5, output t_postbus_type tgt_type_5,
                              input t_postbus_ack tgt_ack_6, output t_postbus_type tgt_type_6,
                              input t_postbus_ack tgt_ack_7, output t_postbus_type tgt_type_7,
                              output t_postbus_data tgt_data
    )
{
    clocked clock rising int_clock reset active_high int_reset t_arb_fsm state = arb_fsm_idle;
    clocked clock rising int_clock reset active_high int_reset bit[3] selected_target = 0 "Target that a current transaction is addressing"; 
    clocked clock rising int_clock reset active_high int_reset bit xfr_first_word = 0 "1 if the source is giving the first word of a transaction";
    comb t_arb_fsm next_state "Next state of FSM";
    comb bit wait "Set if a transfer is in place and the selected target indicates no acknowledge";
    comb t_postbus_type tgt_type "Multiplexed source to target type, which is sent to selected_target if we are active";
    comb t_postbus_ack tgt_ack "Multiplexed target ack, which comes from selected_target if we are active and goes to chosen source";

    /*b Arbitration FSM - state, next_state, wait
     */
    arb_fsm "Arbitration FSM  - select next source to transfer; this is more complex than it need be, as it allows for back-to-back transfers from different masters. But it also does not care about the target of the sources, whereas it could check the target availability for each source first.":
        { 
            next_state = state;
            wait = 0;
            if (state!=arb_fsm_idle)
            {
                wait = (tgt_ack!=0);
            }
            full_switch (state)
                {
                case arb_fsm_idle:
                {   
                    if (src_type_3==postbus_word_type_start) { next_state = arb_fsm_xfr_3; }
                    if (src_type_2==postbus_word_type_start) { next_state = arb_fsm_xfr_2; }
                    if (src_type_1==postbus_word_type_start) { next_state = arb_fsm_xfr_1; }
                    if (src_type_0==postbus_word_type_start) { next_state = arb_fsm_xfr_0; }
                }
                case arb_fsm_xfr_0:
                {
                    if ( (src_type_0==postbus_word_type_last) || ((xfr_first_word) && (src_data_0[0])) )
                    {
                        next_state = arb_fsm_idle;
                        if (src_type_3==postbus_word_type_start) { next_state = arb_fsm_xfr_3; }
                        if (src_type_2==postbus_word_type_start) { next_state = arb_fsm_xfr_2; }
                        if (src_type_1==postbus_word_type_start) { next_state = arb_fsm_xfr_1; }
                    }
                }
                case arb_fsm_xfr_1:
                {
                    if ( (src_type_1==postbus_word_type_last) || ((xfr_first_word) && (src_data_1[0])) )
                    {
                        next_state = arb_fsm_idle;
                        if (src_type_0==postbus_word_type_start) { next_state = arb_fsm_xfr_0; }
                        if (src_type_3==postbus_word_type_start) { next_state = arb_fsm_xfr_3; }
                        if (src_type_2==postbus_word_type_start) { next_state = arb_fsm_xfr_2; }
                    }
                }
                case arb_fsm_xfr_2:
                {
                    if ( (src_type_2==postbus_word_type_last) || ((xfr_first_word) && (src_data_2[0])) )
                    {
                        next_state = arb_fsm_idle;
                        if (src_type_1==postbus_word_type_start) { next_state = arb_fsm_xfr_1; }
                        if (src_type_0==postbus_word_type_start) { next_state = arb_fsm_xfr_0; }
                        if (src_type_3==postbus_word_type_start) { next_state = arb_fsm_xfr_3; }
                    }
                }
                case arb_fsm_xfr_3:
                {
                    if ( (src_type_3==postbus_word_type_last) || ((xfr_first_word) && (src_data_3[0])) )
                    {
                        next_state = arb_fsm_idle;
                        if (src_type_2==postbus_word_type_start) { next_state = arb_fsm_xfr_2; }
                        if (src_type_1==postbus_word_type_start) { next_state = arb_fsm_xfr_1; }
                        if (src_type_0==postbus_word_type_start) { next_state = arb_fsm_xfr_0; }
                    }
                }
                }
            if (wait)
            {
                next_state = state;
            }
            state <= next_state;
        }

    /*b Determine first cycle of a transaction - xfr_first_word
     */
    first_of_transaction "Determine first cycle of a transaction":
        {
            xfr_first_word <= 0;
            if (next_state != state)
            {
                xfr_first_word <= 1;
            }
        }

    /*b Get selected target - selected_target
     */
    select_target "Select target, on change to new target, which is when we change state":
        {
            if (next_state != state)
            {
                full_switch (next_state)
                {
                case arb_fsm_idle:
                case arb_fsm_xfr_0:
                { selected_target <= src_data_0[3;1]; }
                case arb_fsm_xfr_1: {selected_target <= src_data_1[3;1];}
                case arb_fsm_xfr_2: {selected_target <= src_data_2[3;1];}
                case arb_fsm_xfr_3: {selected_target <= src_data_3[3;1];}
                }
            }
        }

    /*b Output muxes for data and target - tgt_data, tgt_type, tgt_type_*, tgt_ack, src_ack_*
     */
    output_mux "Output data, type multiplexers":
        {
            full_switch(state)
                {
                case arb_fsm_idle:
                {
                    tgt_data = src_data_0;
                    tgt_type = postbus_word_type_idle;
                }
                case arb_fsm_xfr_0: 
                {
                    tgt_data = src_data_0;
                    tgt_type = src_type_0;
                }
                case arb_fsm_xfr_1: 
                {
                    tgt_data = src_data_1;
                    tgt_type = src_type_0;
                }
                case arb_fsm_xfr_2: 
                {
                    tgt_data = src_data_2;
                    tgt_type = src_type_0;
                }
                case arb_fsm_xfr_3: 
                {
                    tgt_data = src_data_3;
                    tgt_type = src_type_0;
                }
                }
            tgt_type_0 = postbus_word_type_idle;
            tgt_type_1 = postbus_word_type_idle;
            tgt_type_2 = postbus_word_type_idle;
            tgt_type_3 = postbus_word_type_idle;
            tgt_type_4 = postbus_word_type_idle;
            tgt_type_5 = postbus_word_type_idle;
            tgt_type_6 = postbus_word_type_idle;
            tgt_type_7 = postbus_word_type_idle;
            full_switch( selected_target )
                {
                case 0: {tgt_type_0 = tgt_type; tgt_ack = tgt_ack_0;}
                case 1: {tgt_type_1 = tgt_type; tgt_ack = tgt_ack_1;}
                case 2: {tgt_type_2 = tgt_type; tgt_ack = tgt_ack_2;}
                case 3: {tgt_type_3 = tgt_type; tgt_ack = tgt_ack_3;}
                case 4: {tgt_type_4 = tgt_type; tgt_ack = tgt_ack_4;}
                case 5: {tgt_type_5 = tgt_type; tgt_ack = tgt_ack_5;}
                case 6: {tgt_type_6 = tgt_type; tgt_ack = tgt_ack_6;}
                case 7: {tgt_type_7 = tgt_type; tgt_ack = tgt_ack_7;}
                }

            src_ack_0 = 0;
            src_ack_1 = 0;
            src_ack_2 = 0;
            src_ack_3 = 0;
            part_switch(state)
                {
                case arb_fsm_xfr_0: {src_ack_0 = tgt_ack;}
                case arb_fsm_xfr_1: {src_ack_1 = tgt_ack;}
                case arb_fsm_xfr_2: {src_ack_2 = tgt_ack;}
                case arb_fsm_xfr_3: {src_ack_3 = tgt_ack;}
                }
        }
}
