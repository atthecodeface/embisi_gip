/*a Copyright Gavin J Stark, 2004
 */

/*a To do
 */

/*a Includes
 */
include "io_cmd.h"
include "io_ethernet_rx.h"
include "io_sync_request.h"
include "io_baud_rate_generator.h"
include "io_simple_fifo.h"
include "memories.h"

/*a Constants
 */
constant integer ingress_sram_log_size=9;

/*a Types
 */
/*t t_status_op
 */
typedef enum [2]
{
    status_op_none,
    status_op_write_time,
    status_op_write_data,
} t_status_op;

/*t t_ingress_sram_data_op
 */
typedef enum [2]
{
    ingress_sram_data_op_write_time,
    ingress_sram_data_op_write_status,
    ingress_sram_data_op_write_rx_data,
    ingress_sram_data_op_read
} t_ingress_sram_data_op;

/*t t_ingress_sram_data_reg_op
 */
typedef enum [2]
{
    ingress_sram_data_reg_op_hold,
    ingress_sram_data_reg_op_rx_data,
    ingress_sram_data_reg_op_status,
} t_ingress_sram_data_reg_op;

/*t t_ingress_sram_address_op
 */
typedef enum [2]
{
    ingress_sram_address_op_fifo_read,
    ingress_sram_address_op_fifo_write,
    ingress_sram_address_op_ingress_addressed,
    ingress_sram_address_op_postbus_addressed,
} t_ingress_sram_address_op;

/*a io_block module
 */
module io_block( clock io_clock,
                 input bit io_reset,

                 clock int_clock,
                 input bit int_reset,

                 input bit mii_dv, // goes high during the preamble OR at the latest at the start of the SFD
                 input bit mii_err, // if goes high with dv, then abort the receive; wait until dv goes low
                 input bit[4] mii_data
    )
{
    /*b Variables
     */
    default clock int_clock;
    default reset int_reset;

    net bit[32]               erx_data_fifo_data;
    net t_io_rx_data_fifo_cmd erx_data_fifo_cmd;
    net bit                   erx_data_fifo_toggle;
    net bit                   erx_rxd_req;
    comb bit                   erx_rxd_ack;
    net bit                   erx_data_fifo_full;


    net bit[32]               erx_status_fifo_data;
    net t_io_status_fifo_cmd  erx_status_fifo_cmd;
    net bit                   erx_status_fifo_toggle;
    net bit                   erx_status_req;
    comb bit                   erx_status_ack;

    clocked bit[32] status_timer = 0;
    clocked bit[32] status_data = 0;
    clocked bit status_source = 0;
    clocked t_status_op status_op = status_op_none;

    comb bit ingress_sram_write;
    comb bit ingress_sram_read;
    comb bit[ingress_sram_log_size] ingress_sram_address;
    comb bit[32] ingress_sram_write_data;
    net bit[32] ingress_sram_read_data;

    comb t_simple_fifo_op status_fifo_ptr_op;
    net bit [ingress_sram_log_size-1] status_fifo_write_address;
    net bit [ingress_sram_log_size-1] status_fifo_read_address;
    net bit status_fifo_empty;
    net bit status_fifo_full;
    net bit status_fifo_watermark;
    net bit status_fifo_overflowed;
    net bit status_fifo_underflowed;
    net bit[ingress_sram_log_size-1] cfg_base_address;
    net bit[ingress_sram_log_size-1] cfg_size_m_one;
    net bit[ingress_sram_log_size-1] cfg_watermark;

    comb t_simple_fifo_op rxd_fifo_ptr_op;
    comb bit [ingress_sram_log_size-1] rxd_fifo_write_address;

    net bit brg0_enable;
    comb bit brg0_set_config;
    comb bit[32] config_data;

    /*b Ethernet receive 0 instantiation
     */
    ethernet_receive "Ethernet receive module and sync interface":
        {
            ethernet_rx erx( io_clock <- io_clock,
                             io_reset <= io_reset,

                             data_fifo_data   => erx_data_fifo_data,
                             data_fifo_cmd    => erx_data_fifo_cmd,
                             data_fifo_toggle => erx_data_fifo_toggle,
                             data_fifo_full    = erx_data_fifo_full,

                             status_fifo_data   => erx_status_fifo_data,
                             status_fifo_cmd    => erx_status_fifo_cmd,
                             status_fifo_toggle => erx_status_fifo_toggle,

                             mii_dv <= mii_dv,
                             mii_err <= mii_err,
                             mii_data <= mii_data );

            io_sync_request erx_sr_rxd( int_clock <- int_clock,
                                        int_reset <= int_reset,
                                        io_cmd_toggle <= erx_data_fifo_toggle,
                                        io_arb_request => erx_rxd_req,
                                        arb_io_ack <= erx_rxd_ack );

            io_sync_request erx_sr_status( int_clock <- int_clock,
                                           int_reset <= int_reset,
                                           io_cmd_toggle <= erx_status_fifo_toggle,
                                           io_arb_request => erx_status_req,
                                           arb_io_ack <= erx_status_ack );
        }

    /*b Status and RxData FIFO ptrs and their arbiter
     */
    status_fifos "Status fifos":
        {
            status_timer <= status_timer+1;
            erx_status_ack = 0;
            // Actually we need to take 4 status and 4 rx data requests and a postbus read request, and decide what to do for address calc in cycle+1, with data in cycle+2
            // So postbus requests need to know how many words they want to read; the ack for postbus can be same cycle, though.
            // So we will build a module that takes the 4 status and data requests, returns acks, and pipelined address/data operations (including FIFO number & read/write ptr / address specifier indications)
            // So ingress_sram_op can be:
            //   write timer value
            //   write ingress status data value
            //   write ingress rx data value
            //   ?write postbus data value
            //   read
            // ingress_sram_address can be:
            //   status FIFO 'n' read ptr
            //   status FIFO 'n' write ptr
            //   postbus address
            //   ingress status address value
            // data reg op can be
            //   hold
            //   record ingress rx data port 'n'
            //   record ingress status port 'n'
            // address reg op can be
            //   hold
            //   record ingress rx data address 'n' (status is always FIFO)
            full_switch( status_op )
                {
                case status_op_none:
                {
                    if (erx_status_req)
                    {
                        status_op <= status_op_write_time;
                        status_data <= erx_status_fifo_data;
                    }
                }
                case status_op_write_time:
                {
                    status_op <= status_op_write_data;
                    erx_status_ack = 1;
                    ingress_sram_write = 1;
                    ingress_sram_write_data = status_timer;
                    ingress_sram_address[ingress_sram_log_size-1;1] = status_fifo_write_address;
                    ingress_sram_address[0] = 0;
                }
                case status_op_write_data: // also arbitrate for next user; unless a data is pending, in which case go to none anyway so data can be written (interleave status and data writes)
                {
                    status_op <= status_op_none;
                    status_fifo_ptr_op = simple_fifo_op_inc_write_ptr;
                    ingress_sram_write = 1;
                    ingress_sram_write_data = status_data;
                    ingress_sram_address[ingress_sram_log_size-1;1] = status_fifo_write_address;
                    ingress_sram_address[0] = 1;
                }
                }
            io_simple_fifo status_fifo_ptrs( int_clock <- int_clock,
                                             int_reset <= int_reset,
                                             fifo_op <= status_fifo_ptr_op,
                                             fifo_write_address => status_fifo_write_address,
                                             fifo_read_address => status_fifo_read_address,
                                             fifo_empty => status_fifo_empty,
                                             fifo_full => status_fifo_full,
                                             fifo_watermark => status_fifo_watermark,
                                             fifo_overflowed => status_fifo_overflowed,
                                             fifo_underflowed => status_fifo_underflowed,
                                             cfg_base_address <= cfg_base_address,
                                             cfg_size_m_one <= cfg_size_m_one,
                                             cfg_watermark <= cfg_watermark );

        }

    /*b Ingress SRAM operation, data and address selectors
     */
    status_fifos "Status fifos":
        {
            /*b Status timer
             */
            status_timer <= status_timer+1;

            /*b Handle the data op
             */
            //   write timer value
            //   write ingress status data value
            //   write ingress rx data value
            //   ?write postbus data value
            //   read
            ingress_sram_write = 0;
            ingress_sram_read = 0;
            ingress_sram_write_data = ingress_data_reg;
            full_switch ( ingress_sram_data_op )
                {
                case ingress_sram_data_op_write_time:
                {
                    ingress_sram_write = 1;
                    ingress_sram_write_data = status_timer;
                }
                case ingress_sram_data_op_write_status:
                case ingress_sram_data_op_write_rx_data:
                {
                    ingress_sram_write = 1;
                    ingress_sram_write_data = ingress_data_reg;
                }
                case ingress_sram_data_op_read:
                {
                    ingress_sram_read = 1;
                    ingress_sram_write_data = ingress_data_reg;
                }
                }

            /*b Handle the data reg - should select the appropriate interface, but we have just one at present
             */
            full_switch ( ingress_sram_data_reg_op )
                {
                case ingress_sram_data_reg_op_hold:
                {
                }
                case ingress_sram_data_reg_op_rx_data:
                {
                    ingress_data_reg <= erx_data_fifo_data;
                }
                case ingress_sram_data_reg_op_status:
                {
                    ingress_data_reg <= erx_status_fifo_data;
                }
                }

            /*b Handle the SRAM address
             */
            full_switch ( ingress_sram_address_op )
                {
                case ingress_sram_address_op_fifo_read:
                case ingress_sram_address_op_fifo_write:
                {
                    ingress_sram_address = ingress_fifo_address;
                }
                case ingress_sram_address_op_ingress_addressed:
                {
                    //ingress_sram_address = ingress_data_address;
                }
                case ingress_sram_address_op_postbus_addressed:
                {
                    //ingress_sram_address = ingress_postbus_address;
                }
        }

    /*b Ingress SRAM (RxDatat and status)
     */
    ingress_sram "Ingress sram":
        {
            memory_s_sp_2048_x_32 ingress_sram( sram_clock <- int_clock,
                                                sram_read <= ingress_sram_read,
                                                sram_write <= ingress_sram_write,
                                                sram_address <= ingress_sram_address,
                                                sram_write_data <= ingress_sram_write_data,
                                                sram_read_data => ingress_sram_read_data );
        }

    /*b Baud rate generators
     */
    brg "Baud rate generators":
        {
            io_baud_rate_generator brg0 ( io_clock <- io_clock,
                                          io_reset <= io_reset,
                                          counter_enable <= 1, // or allow for daisychaining or divide-by-input-enable
                                          counter_reset <= 0, // or allow for synchronization
                                          baud_clock_enable => brg0_enable,
                                          set_clock_config <= brg0_set_config,
                                          config_baud_addition_value <= config_data[io_baud_rate_divider_size;0], // Bottom sixteen bits contain the addition value
                                          config_baud_subtraction_value <= config_data[io_baud_rate_divider_size;16] // Top sixteen bits contain the addition value
                );
        }

    /*b Done
     */
}
