/*a Copyright Gavin J Stark, 2004
 */

/*a To do
 */

/*a Includes
 */
include "io_sync_request.h"

/*a Constants
 */

/*a Types
 */
typedef struct
{
    bit[2] regs;
    bit value;
} t_sync;

/*a io_sync_request module
 */
module io_sync_request(
	 clock int_clock "main system clck",
	 input bit int_reset "main system reset",
	 input bit io_cmd_toggle "Toggle from IO clock domain that indicates a request",
	 output bit io_arb_request "Actual request to arbiter, derived directly from registers",
	 input bit arb_io_ack "Combinatorial acknowledge of request" )
	"This module synchronizes a request for a command execution and requests that of the arbiter, removing the request when it has been acknowledged"
{
	 default clock int_clock;
	 default reset int_reset;

     clocked t_sync sync = { regs=0, value=0 } "Synchronizer for the toggle";
	 clocked bit request_pending=0;

	 comb bit request_just_arrived;

     sync_and_req "Synchronizers and request":
         {
             sync.regs[0] <= io_cmd_toggle;
             sync.regs[1] <= sync.regs[0];
             sync.value <= sync.regs[1];
             request_just_arrived = (sync.value != sync.regs[1]);
         }

     request_pending "Request pending and out, handling acknowledge":
         {
             if (arb_io_ack)
             {
                 request_pending <= 0;
             }
             elsif (request_just_arrived)
                 {
                     request_pending <= 1;
                 }

             io_arb_request = 0;
             if ( request_just_arrived || request_pending )
             {
                 io_arb_request = 1;
             }
         }
}
