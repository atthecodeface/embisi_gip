module barrel_shift_32
(
    select, in, out
);
input [4:0]select;
input [31:0]in;
output [31:0]out;
wire [31:0] stage_1;
wire [31:0] stage_2;
wire [31:0] stage_3;
wire [31:0] stage_4;
wire [31:0] stage_5;

    // A MUX is a LUT3 where the inputs / output are as follows
    // I2==S  I1  I0   O
    //     0   0   0   0
    //     0   0   1   1
    //     0   1   0   0
    //     0   1   1   1
    //     1   0   0   0
    //     1   0   1   0
    //     1   1   0   1
    //     1   1   1   1
    // So the LUT3 init is ca

    LUT3 mux_1_00 ( .O(stage_1[ 0]), .I0( in[ 0] ), .I1( in[16] ), .I2( select[4] ) ); defparam mux_1_00.INIT = 8'hca; //'
    LUT3 mux_1_01 ( .O(stage_1[ 1]), .I0( in[ 1] ), .I1( in[17] ), .I2( select[4] ) ); defparam mux_1_01.INIT = 8'hca; //'
    LUT3 mux_1_02 ( .O(stage_1[ 2]), .I0( in[ 2] ), .I1( in[18] ), .I2( select[4] ) ); defparam mux_1_02.INIT = 8'hca; //'
    LUT3 mux_1_03 ( .O(stage_1[ 3]), .I0( in[ 3] ), .I1( in[19] ), .I2( select[4] ) ); defparam mux_1_03.INIT = 8'hca; //'
    LUT3 mux_1_04 ( .O(stage_1[ 4]), .I0( in[ 4] ), .I1( in[20] ), .I2( select[4] ) ); defparam mux_1_04.INIT = 8'hca; //'
    LUT3 mux_1_05 ( .O(stage_1[ 5]), .I0( in[ 5] ), .I1( in[21] ), .I2( select[4] ) ); defparam mux_1_05.INIT = 8'hca; //'
    LUT3 mux_1_06 ( .O(stage_1[ 6]), .I0( in[ 6] ), .I1( in[22] ), .I2( select[4] ) ); defparam mux_1_06.INIT = 8'hca; //'
    LUT3 mux_1_07 ( .O(stage_1[ 7]), .I0( in[ 7] ), .I1( in[23] ), .I2( select[4] ) ); defparam mux_1_07.INIT = 8'hca; //'
    LUT3 mux_1_08 ( .O(stage_1[ 8]), .I0( in[ 8] ), .I1( in[24] ), .I2( select[4] ) ); defparam mux_1_08.INIT = 8'hca; //'
    LUT3 mux_1_09 ( .O(stage_1[ 9]), .I0( in[ 9] ), .I1( in[25] ), .I2( select[4] ) ); defparam mux_1_09.INIT = 8'hca; //'
    LUT3 mux_1_10 ( .O(stage_1[10]), .I0( in[10] ), .I1( in[26] ), .I2( select[4] ) ); defparam mux_1_10.INIT = 8'hca; //'
    LUT3 mux_1_11 ( .O(stage_1[11]), .I0( in[11] ), .I1( in[27] ), .I2( select[4] ) ); defparam mux_1_11.INIT = 8'hca; //'
    LUT3 mux_1_12 ( .O(stage_1[12]), .I0( in[12] ), .I1( in[28] ), .I2( select[4] ) ); defparam mux_1_12.INIT = 8'hca; //'
    LUT3 mux_1_13 ( .O(stage_1[13]), .I0( in[13] ), .I1( in[29] ), .I2( select[4] ) ); defparam mux_1_13.INIT = 8'hca; //'
    LUT3 mux_1_14 ( .O(stage_1[14]), .I0( in[14] ), .I1( in[30] ), .I2( select[4] ) ); defparam mux_1_14.INIT = 8'hca; //'
    LUT3 mux_1_15 ( .O(stage_1[15]), .I0( in[15] ), .I1( in[31] ), .I2( select[4] ) ); defparam mux_1_15.INIT = 8'hca; //'
    LUT3 mux_1_16 ( .O(stage_1[16]), .I0( in[16] ), .I1( in[ 0] ), .I2( select[4] ) ); defparam mux_1_16.INIT = 8'hca; //'
    LUT3 mux_1_17 ( .O(stage_1[17]), .I0( in[17] ), .I1( in[ 1] ), .I2( select[4] ) ); defparam mux_1_17.INIT = 8'hca; //'
    LUT3 mux_1_18 ( .O(stage_1[18]), .I0( in[18] ), .I1( in[ 2] ), .I2( select[4] ) ); defparam mux_1_18.INIT = 8'hca; //'
    LUT3 mux_1_19 ( .O(stage_1[19]), .I0( in[19] ), .I1( in[ 3] ), .I2( select[4] ) ); defparam mux_1_19.INIT = 8'hca; //'
    LUT3 mux_1_20 ( .O(stage_1[20]), .I0( in[20] ), .I1( in[ 4] ), .I2( select[4] ) ); defparam mux_1_20.INIT = 8'hca; //'
    LUT3 mux_1_21 ( .O(stage_1[21]), .I0( in[21] ), .I1( in[ 5] ), .I2( select[4] ) ); defparam mux_1_21.INIT = 8'hca; //'
    LUT3 mux_1_22 ( .O(stage_1[22]), .I0( in[22] ), .I1( in[ 6] ), .I2( select[4] ) ); defparam mux_1_22.INIT = 8'hca; //'
    LUT3 mux_1_23 ( .O(stage_1[23]), .I0( in[23] ), .I1( in[ 7] ), .I2( select[4] ) ); defparam mux_1_23.INIT = 8'hca; //'
    LUT3 mux_1_24 ( .O(stage_1[24]), .I0( in[24] ), .I1( in[ 8] ), .I2( select[4] ) ); defparam mux_1_24.INIT = 8'hca; //'
    LUT3 mux_1_25 ( .O(stage_1[25]), .I0( in[25] ), .I1( in[ 9] ), .I2( select[4] ) ); defparam mux_1_25.INIT = 8'hca; //'
    LUT3 mux_1_26 ( .O(stage_1[26]), .I0( in[26] ), .I1( in[10] ), .I2( select[4] ) ); defparam mux_1_26.INIT = 8'hca; //'
    LUT3 mux_1_27 ( .O(stage_1[27]), .I0( in[27] ), .I1( in[11] ), .I2( select[4] ) ); defparam mux_1_27.INIT = 8'hca; //'
    LUT3 mux_1_28 ( .O(stage_1[28]), .I0( in[28] ), .I1( in[12] ), .I2( select[4] ) ); defparam mux_1_28.INIT = 8'hca; //'
    LUT3 mux_1_29 ( .O(stage_1[29]), .I0( in[29] ), .I1( in[13] ), .I2( select[4] ) ); defparam mux_1_29.INIT = 8'hca; //'
    LUT3 mux_1_30 ( .O(stage_1[30]), .I0( in[30] ), .I1( in[14] ), .I2( select[4] ) ); defparam mux_1_30.INIT = 8'hca; //'
    LUT3 mux_1_31 ( .O(stage_1[31]), .I0( in[31] ), .I1( in[15] ), .I2( select[4] ) ); defparam mux_1_31.INIT = 8'hca; //'

    LUT3 mux_2_00 ( .O(stage_2[ 0]), .I0( stage_1[ 0] ), .I1( stage_1[ 8] ), .I2( select[3] ) ); defparam mux_2_00.INIT = 8'hca; //'
    LUT3 mux_2_01 ( .O(stage_2[ 1]), .I0( stage_1[ 1] ), .I1( stage_1[ 9] ), .I2( select[3] ) ); defparam mux_2_01.INIT = 8'hca; //'
    LUT3 mux_2_02 ( .O(stage_2[ 2]), .I0( stage_1[ 2] ), .I1( stage_1[10] ), .I2( select[3] ) ); defparam mux_2_02.INIT = 8'hca; //'
    LUT3 mux_2_03 ( .O(stage_2[ 3]), .I0( stage_1[ 3] ), .I1( stage_1[11] ), .I2( select[3] ) ); defparam mux_2_03.INIT = 8'hca; //'
    LUT3 mux_2_04 ( .O(stage_2[ 4]), .I0( stage_1[ 4] ), .I1( stage_1[12] ), .I2( select[3] ) ); defparam mux_2_04.INIT = 8'hca; //'
    LUT3 mux_2_05 ( .O(stage_2[ 5]), .I0( stage_1[ 5] ), .I1( stage_1[13] ), .I2( select[3] ) ); defparam mux_2_05.INIT = 8'hca; //'
    LUT3 mux_2_06 ( .O(stage_2[ 6]), .I0( stage_1[ 6] ), .I1( stage_1[14] ), .I2( select[3] ) ); defparam mux_2_06.INIT = 8'hca; //'
    LUT3 mux_2_07 ( .O(stage_2[ 7]), .I0( stage_1[ 7] ), .I1( stage_1[15] ), .I2( select[3] ) ); defparam mux_2_07.INIT = 8'hca; //'
    LUT3 mux_2_08 ( .O(stage_2[ 8]), .I0( stage_1[ 8] ), .I1( stage_1[16] ), .I2( select[3] ) ); defparam mux_2_08.INIT = 8'hca; //'
    LUT3 mux_2_09 ( .O(stage_2[ 9]), .I0( stage_1[ 9] ), .I1( stage_1[17] ), .I2( select[3] ) ); defparam mux_2_09.INIT = 8'hca; //'
    LUT3 mux_2_10 ( .O(stage_2[10]), .I0( stage_1[10] ), .I1( stage_1[18] ), .I2( select[3] ) ); defparam mux_2_10.INIT = 8'hca; //'
    LUT3 mux_2_11 ( .O(stage_2[11]), .I0( stage_1[11] ), .I1( stage_1[19] ), .I2( select[3] ) ); defparam mux_2_11.INIT = 8'hca; //'
    LUT3 mux_2_12 ( .O(stage_2[12]), .I0( stage_1[12] ), .I1( stage_1[20] ), .I2( select[3] ) ); defparam mux_2_12.INIT = 8'hca; //'
    LUT3 mux_2_13 ( .O(stage_2[13]), .I0( stage_1[13] ), .I1( stage_1[21] ), .I2( select[3] ) ); defparam mux_2_13.INIT = 8'hca; //'
    LUT3 mux_2_14 ( .O(stage_2[14]), .I0( stage_1[14] ), .I1( stage_1[22] ), .I2( select[3] ) ); defparam mux_2_14.INIT = 8'hca; //'
    LUT3 mux_2_15 ( .O(stage_2[15]), .I0( stage_1[15] ), .I1( stage_1[23] ), .I2( select[3] ) ); defparam mux_2_15.INIT = 8'hca; //'
    LUT3 mux_2_16 ( .O(stage_2[16]), .I0( stage_1[16] ), .I1( stage_1[24] ), .I2( select[3] ) ); defparam mux_2_16.INIT = 8'hca; //'
    LUT3 mux_2_17 ( .O(stage_2[17]), .I0( stage_1[17] ), .I1( stage_1[25] ), .I2( select[3] ) ); defparam mux_2_17.INIT = 8'hca; //'
    LUT3 mux_2_18 ( .O(stage_2[18]), .I0( stage_1[18] ), .I1( stage_1[26] ), .I2( select[3] ) ); defparam mux_2_18.INIT = 8'hca; //'
    LUT3 mux_2_19 ( .O(stage_2[19]), .I0( stage_1[19] ), .I1( stage_1[27] ), .I2( select[3] ) ); defparam mux_2_19.INIT = 8'hca; //'
    LUT3 mux_2_20 ( .O(stage_2[20]), .I0( stage_1[20] ), .I1( stage_1[28] ), .I2( select[3] ) ); defparam mux_2_20.INIT = 8'hca; //'
    LUT3 mux_2_21 ( .O(stage_2[21]), .I0( stage_1[21] ), .I1( stage_1[29] ), .I2( select[3] ) ); defparam mux_2_21.INIT = 8'hca; //'
    LUT3 mux_2_22 ( .O(stage_2[22]), .I0( stage_1[22] ), .I1( stage_1[30] ), .I2( select[3] ) ); defparam mux_2_22.INIT = 8'hca; //'
    LUT3 mux_2_23 ( .O(stage_2[23]), .I0( stage_1[23] ), .I1( stage_1[31] ), .I2( select[3] ) ); defparam mux_2_23.INIT = 8'hca; //'
    LUT3 mux_2_24 ( .O(stage_2[24]), .I0( stage_1[24] ), .I1( stage_1[ 0] ), .I2( select[3] ) ); defparam mux_2_24.INIT = 8'hca; //'
    LUT3 mux_2_25 ( .O(stage_2[25]), .I0( stage_1[25] ), .I1( stage_1[ 1] ), .I2( select[3] ) ); defparam mux_2_25.INIT = 8'hca; //'
    LUT3 mux_2_26 ( .O(stage_2[26]), .I0( stage_1[26] ), .I1( stage_1[ 2] ), .I2( select[3] ) ); defparam mux_2_26.INIT = 8'hca; //'
    LUT3 mux_2_27 ( .O(stage_2[27]), .I0( stage_1[27] ), .I1( stage_1[ 3] ), .I2( select[3] ) ); defparam mux_2_27.INIT = 8'hca; //'
    LUT3 mux_2_28 ( .O(stage_2[28]), .I0( stage_1[28] ), .I1( stage_1[ 4] ), .I2( select[3] ) ); defparam mux_2_28.INIT = 8'hca; //'
    LUT3 mux_2_29 ( .O(stage_2[29]), .I0( stage_1[29] ), .I1( stage_1[ 5] ), .I2( select[3] ) ); defparam mux_2_29.INIT = 8'hca; //'
    LUT3 mux_2_30 ( .O(stage_2[30]), .I0( stage_1[30] ), .I1( stage_1[ 6] ), .I2( select[3] ) ); defparam mux_2_30.INIT = 8'hca; //'
    LUT3 mux_2_31 ( .O(stage_2[31]), .I0( stage_1[31] ), .I1( stage_1[ 7] ), .I2( select[3] ) ); defparam mux_2_31.INIT = 8'hca; //'

    LUT3 mux_3_00 ( .O(stage_3[ 0]), .I0( stage_2[ 0] ), .I1( stage_2[ 4] ), .I2( select[2] ) ); defparam mux_3_00.INIT = 8'hca; //'
    LUT3 mux_3_01 ( .O(stage_3[ 1]), .I0( stage_2[ 1] ), .I1( stage_2[ 5] ), .I2( select[2] ) ); defparam mux_3_01.INIT = 8'hca; //'
    LUT3 mux_3_02 ( .O(stage_3[ 2]), .I0( stage_2[ 2] ), .I1( stage_2[ 6] ), .I2( select[2] ) ); defparam mux_3_02.INIT = 8'hca; //'
    LUT3 mux_3_03 ( .O(stage_3[ 3]), .I0( stage_2[ 3] ), .I1( stage_2[ 7] ), .I2( select[2] ) ); defparam mux_3_03.INIT = 8'hca; //'
    LUT3 mux_3_04 ( .O(stage_3[ 4]), .I0( stage_2[ 4] ), .I1( stage_2[ 8] ), .I2( select[2] ) ); defparam mux_3_04.INIT = 8'hca; //'
    LUT3 mux_3_05 ( .O(stage_3[ 5]), .I0( stage_2[ 5] ), .I1( stage_2[ 9] ), .I2( select[2] ) ); defparam mux_3_05.INIT = 8'hca; //'
    LUT3 mux_3_06 ( .O(stage_3[ 6]), .I0( stage_2[ 6] ), .I1( stage_2[10] ), .I2( select[2] ) ); defparam mux_3_06.INIT = 8'hca; //'
    LUT3 mux_3_07 ( .O(stage_3[ 7]), .I0( stage_2[ 7] ), .I1( stage_2[11] ), .I2( select[2] ) ); defparam mux_3_07.INIT = 8'hca; //'
    LUT3 mux_3_08 ( .O(stage_3[ 8]), .I0( stage_2[ 8] ), .I1( stage_2[12] ), .I2( select[2] ) ); defparam mux_3_08.INIT = 8'hca; //'
    LUT3 mux_3_09 ( .O(stage_3[ 9]), .I0( stage_2[ 9] ), .I1( stage_2[13] ), .I2( select[2] ) ); defparam mux_3_09.INIT = 8'hca; //'
    LUT3 mux_3_10 ( .O(stage_3[10]), .I0( stage_2[10] ), .I1( stage_2[14] ), .I2( select[2] ) ); defparam mux_3_10.INIT = 8'hca; //'
    LUT3 mux_3_11 ( .O(stage_3[11]), .I0( stage_2[11] ), .I1( stage_2[15] ), .I2( select[2] ) ); defparam mux_3_11.INIT = 8'hca; //'
    LUT3 mux_3_12 ( .O(stage_3[12]), .I0( stage_2[12] ), .I1( stage_2[16] ), .I2( select[2] ) ); defparam mux_3_12.INIT = 8'hca; //'
    LUT3 mux_3_13 ( .O(stage_3[13]), .I0( stage_2[13] ), .I1( stage_2[17] ), .I2( select[2] ) ); defparam mux_3_13.INIT = 8'hca; //'
    LUT3 mux_3_14 ( .O(stage_3[14]), .I0( stage_2[14] ), .I1( stage_2[18] ), .I2( select[2] ) ); defparam mux_3_14.INIT = 8'hca; //'
    LUT3 mux_3_15 ( .O(stage_3[15]), .I0( stage_2[15] ), .I1( stage_2[19] ), .I2( select[2] ) ); defparam mux_3_15.INIT = 8'hca; //'
    LUT3 mux_3_16 ( .O(stage_3[16]), .I0( stage_2[16] ), .I1( stage_2[20] ), .I2( select[2] ) ); defparam mux_3_16.INIT = 8'hca; //'
    LUT3 mux_3_17 ( .O(stage_3[17]), .I0( stage_2[17] ), .I1( stage_2[21] ), .I2( select[2] ) ); defparam mux_3_17.INIT = 8'hca; //'
    LUT3 mux_3_18 ( .O(stage_3[18]), .I0( stage_2[18] ), .I1( stage_2[22] ), .I2( select[2] ) ); defparam mux_3_18.INIT = 8'hca; //'
    LUT3 mux_3_19 ( .O(stage_3[19]), .I0( stage_2[19] ), .I1( stage_2[23] ), .I2( select[2] ) ); defparam mux_3_19.INIT = 8'hca; //'
    LUT3 mux_3_20 ( .O(stage_3[20]), .I0( stage_2[20] ), .I1( stage_2[24] ), .I2( select[2] ) ); defparam mux_3_20.INIT = 8'hca; //'
    LUT3 mux_3_21 ( .O(stage_3[21]), .I0( stage_2[21] ), .I1( stage_2[25] ), .I2( select[2] ) ); defparam mux_3_21.INIT = 8'hca; //'
    LUT3 mux_3_22 ( .O(stage_3[22]), .I0( stage_2[22] ), .I1( stage_2[26] ), .I2( select[2] ) ); defparam mux_3_22.INIT = 8'hca; //'
    LUT3 mux_3_23 ( .O(stage_3[23]), .I0( stage_2[23] ), .I1( stage_2[27] ), .I2( select[2] ) ); defparam mux_3_23.INIT = 8'hca; //'
    LUT3 mux_3_24 ( .O(stage_3[24]), .I0( stage_2[24] ), .I1( stage_2[28] ), .I2( select[2] ) ); defparam mux_3_24.INIT = 8'hca; //'
    LUT3 mux_3_25 ( .O(stage_3[25]), .I0( stage_2[25] ), .I1( stage_2[29] ), .I2( select[2] ) ); defparam mux_3_25.INIT = 8'hca; //'
    LUT3 mux_3_26 ( .O(stage_3[26]), .I0( stage_2[26] ), .I1( stage_2[30] ), .I2( select[2] ) ); defparam mux_3_26.INIT = 8'hca; //'
    LUT3 mux_3_27 ( .O(stage_3[27]), .I0( stage_2[27] ), .I1( stage_2[31] ), .I2( select[2] ) ); defparam mux_3_27.INIT = 8'hca; //'
    LUT3 mux_3_28 ( .O(stage_3[28]), .I0( stage_2[28] ), .I1( stage_2[ 0] ), .I2( select[2] ) ); defparam mux_3_28.INIT = 8'hca; //'
    LUT3 mux_3_29 ( .O(stage_3[29]), .I0( stage_2[29] ), .I1( stage_2[ 1] ), .I2( select[2] ) ); defparam mux_3_29.INIT = 8'hca; //'
    LUT3 mux_3_30 ( .O(stage_3[30]), .I0( stage_2[30] ), .I1( stage_2[ 2] ), .I2( select[2] ) ); defparam mux_3_30.INIT = 8'hca; //'
    LUT3 mux_3_31 ( .O(stage_3[31]), .I0( stage_2[31] ), .I1( stage_2[ 3] ), .I2( select[2] ) ); defparam mux_3_31.INIT = 8'hca; //'

    LUT3 mux_4_00 ( .O(stage_4[ 0]), .I0( stage_3[ 0] ), .I1( stage_3[ 2] ), .I2( select[1] ) ); defparam mux_4_00.INIT = 8'hca; //'
    LUT3 mux_4_01 ( .O(stage_4[ 1]), .I0( stage_3[ 1] ), .I1( stage_3[ 3] ), .I2( select[1] ) ); defparam mux_4_01.INIT = 8'hca; //'
    LUT3 mux_4_02 ( .O(stage_4[ 2]), .I0( stage_3[ 2] ), .I1( stage_3[ 4] ), .I2( select[1] ) ); defparam mux_4_02.INIT = 8'hca; //'
    LUT3 mux_4_03 ( .O(stage_4[ 3]), .I0( stage_3[ 3] ), .I1( stage_3[ 5] ), .I2( select[1] ) ); defparam mux_4_03.INIT = 8'hca; //'
    LUT3 mux_4_04 ( .O(stage_4[ 4]), .I0( stage_3[ 4] ), .I1( stage_3[ 6] ), .I2( select[1] ) ); defparam mux_4_04.INIT = 8'hca; //'
    LUT3 mux_4_05 ( .O(stage_4[ 5]), .I0( stage_3[ 5] ), .I1( stage_3[ 7] ), .I2( select[1] ) ); defparam mux_4_05.INIT = 8'hca; //'
    LUT3 mux_4_06 ( .O(stage_4[ 6]), .I0( stage_3[ 6] ), .I1( stage_3[ 8] ), .I2( select[1] ) ); defparam mux_4_06.INIT = 8'hca; //'
    LUT3 mux_4_07 ( .O(stage_4[ 7]), .I0( stage_3[ 7] ), .I1( stage_3[ 9] ), .I2( select[1] ) ); defparam mux_4_07.INIT = 8'hca; //'
    LUT3 mux_4_08 ( .O(stage_4[ 8]), .I0( stage_3[ 8] ), .I1( stage_3[10] ), .I2( select[1] ) ); defparam mux_4_08.INIT = 8'hca; //'
    LUT3 mux_4_09 ( .O(stage_4[ 9]), .I0( stage_3[ 9] ), .I1( stage_3[11] ), .I2( select[1] ) ); defparam mux_4_09.INIT = 8'hca; //'
    LUT3 mux_4_10 ( .O(stage_4[10]), .I0( stage_3[10] ), .I1( stage_3[12] ), .I2( select[1] ) ); defparam mux_4_10.INIT = 8'hca; //'
    LUT3 mux_4_11 ( .O(stage_4[11]), .I0( stage_3[11] ), .I1( stage_3[13] ), .I2( select[1] ) ); defparam mux_4_11.INIT = 8'hca; //'
    LUT3 mux_4_12 ( .O(stage_4[12]), .I0( stage_3[12] ), .I1( stage_3[14] ), .I2( select[1] ) ); defparam mux_4_12.INIT = 8'hca; //'
    LUT3 mux_4_13 ( .O(stage_4[13]), .I0( stage_3[13] ), .I1( stage_3[15] ), .I2( select[1] ) ); defparam mux_4_13.INIT = 8'hca; //'
    LUT3 mux_4_14 ( .O(stage_4[14]), .I0( stage_3[14] ), .I1( stage_3[16] ), .I2( select[1] ) ); defparam mux_4_14.INIT = 8'hca; //'
    LUT3 mux_4_15 ( .O(stage_4[15]), .I0( stage_3[15] ), .I1( stage_3[17] ), .I2( select[1] ) ); defparam mux_4_15.INIT = 8'hca; //'
    LUT3 mux_4_16 ( .O(stage_4[16]), .I0( stage_3[16] ), .I1( stage_3[18] ), .I2( select[1] ) ); defparam mux_4_16.INIT = 8'hca; //'
    LUT3 mux_4_17 ( .O(stage_4[17]), .I0( stage_3[17] ), .I1( stage_3[19] ), .I2( select[1] ) ); defparam mux_4_17.INIT = 8'hca; //'
    LUT3 mux_4_18 ( .O(stage_4[18]), .I0( stage_3[18] ), .I1( stage_3[20] ), .I2( select[1] ) ); defparam mux_4_18.INIT = 8'hca; //'
    LUT3 mux_4_19 ( .O(stage_4[19]), .I0( stage_3[19] ), .I1( stage_3[21] ), .I2( select[1] ) ); defparam mux_4_19.INIT = 8'hca; //'
    LUT3 mux_4_20 ( .O(stage_4[20]), .I0( stage_3[20] ), .I1( stage_3[22] ), .I2( select[1] ) ); defparam mux_4_20.INIT = 8'hca; //'
    LUT3 mux_4_21 ( .O(stage_4[21]), .I0( stage_3[21] ), .I1( stage_3[23] ), .I2( select[1] ) ); defparam mux_4_21.INIT = 8'hca; //'
    LUT3 mux_4_22 ( .O(stage_4[22]), .I0( stage_3[22] ), .I1( stage_3[24] ), .I2( select[1] ) ); defparam mux_4_22.INIT = 8'hca; //'
    LUT3 mux_4_23 ( .O(stage_4[23]), .I0( stage_3[23] ), .I1( stage_3[25] ), .I2( select[1] ) ); defparam mux_4_23.INIT = 8'hca; //'
    LUT3 mux_4_24 ( .O(stage_4[24]), .I0( stage_3[24] ), .I1( stage_3[26] ), .I2( select[1] ) ); defparam mux_4_24.INIT = 8'hca; //'
    LUT3 mux_4_25 ( .O(stage_4[25]), .I0( stage_3[25] ), .I1( stage_3[27] ), .I2( select[1] ) ); defparam mux_4_25.INIT = 8'hca; //'
    LUT3 mux_4_26 ( .O(stage_4[26]), .I0( stage_3[26] ), .I1( stage_3[28] ), .I2( select[1] ) ); defparam mux_4_26.INIT = 8'hca; //'
    LUT3 mux_4_27 ( .O(stage_4[27]), .I0( stage_3[27] ), .I1( stage_3[29] ), .I2( select[1] ) ); defparam mux_4_27.INIT = 8'hca; //'
    LUT3 mux_4_28 ( .O(stage_4[28]), .I0( stage_3[28] ), .I1( stage_3[30] ), .I2( select[1] ) ); defparam mux_4_28.INIT = 8'hca; //'
    LUT3 mux_4_29 ( .O(stage_4[29]), .I0( stage_3[29] ), .I1( stage_3[31] ), .I2( select[1] ) ); defparam mux_4_29.INIT = 8'hca; //'
    LUT3 mux_4_30 ( .O(stage_4[30]), .I0( stage_3[30] ), .I1( stage_3[ 0] ), .I2( select[1] ) ); defparam mux_4_30.INIT = 8'hca; //'
    LUT3 mux_4_31 ( .O(stage_4[31]), .I0( stage_3[31] ), .I1( stage_3[ 1] ), .I2( select[1] ) ); defparam mux_4_31.INIT = 8'hca; //'

    LUT3 mux_5_00 ( .O(stage_5[ 0]), .I0( stage_4[ 0] ), .I1( stage_4[ 1] ), .I2( select[0] ) ); defparam mux_5_00.INIT = 8'hca; //'
    LUT3 mux_5_01 ( .O(stage_5[ 1]), .I0( stage_4[ 1] ), .I1( stage_4[ 2] ), .I2( select[0] ) ); defparam mux_5_01.INIT = 8'hca; //'
    LUT3 mux_5_02 ( .O(stage_5[ 2]), .I0( stage_4[ 2] ), .I1( stage_4[ 3] ), .I2( select[0] ) ); defparam mux_5_02.INIT = 8'hca; //'
    LUT3 mux_5_03 ( .O(stage_5[ 3]), .I0( stage_4[ 3] ), .I1( stage_4[ 4] ), .I2( select[0] ) ); defparam mux_5_03.INIT = 8'hca; //'
    LUT3 mux_5_04 ( .O(stage_5[ 4]), .I0( stage_4[ 4] ), .I1( stage_4[ 5] ), .I2( select[0] ) ); defparam mux_5_04.INIT = 8'hca; //'
    LUT3 mux_5_05 ( .O(stage_5[ 5]), .I0( stage_4[ 5] ), .I1( stage_4[ 6] ), .I2( select[0] ) ); defparam mux_5_05.INIT = 8'hca; //'
    LUT3 mux_5_06 ( .O(stage_5[ 6]), .I0( stage_4[ 6] ), .I1( stage_4[ 7] ), .I2( select[0] ) ); defparam mux_5_06.INIT = 8'hca; //'
    LUT3 mux_5_07 ( .O(stage_5[ 7]), .I0( stage_4[ 7] ), .I1( stage_4[ 8] ), .I2( select[0] ) ); defparam mux_5_07.INIT = 8'hca; //'
    LUT3 mux_5_08 ( .O(stage_5[ 8]), .I0( stage_4[ 8] ), .I1( stage_4[ 9] ), .I2( select[0] ) ); defparam mux_5_08.INIT = 8'hca; //'
    LUT3 mux_5_09 ( .O(stage_5[ 9]), .I0( stage_4[ 9] ), .I1( stage_4[10] ), .I2( select[0] ) ); defparam mux_5_09.INIT = 8'hca; //'
    LUT3 mux_5_10 ( .O(stage_5[10]), .I0( stage_4[10] ), .I1( stage_4[11] ), .I2( select[0] ) ); defparam mux_5_10.INIT = 8'hca; //'
    LUT3 mux_5_11 ( .O(stage_5[11]), .I0( stage_4[11] ), .I1( stage_4[12] ), .I2( select[0] ) ); defparam mux_5_11.INIT = 8'hca; //'
    LUT3 mux_5_12 ( .O(stage_5[12]), .I0( stage_4[12] ), .I1( stage_4[13] ), .I2( select[0] ) ); defparam mux_5_12.INIT = 8'hca; //'
    LUT3 mux_5_13 ( .O(stage_5[13]), .I0( stage_4[13] ), .I1( stage_4[14] ), .I2( select[0] ) ); defparam mux_5_13.INIT = 8'hca; //'
    LUT3 mux_5_14 ( .O(stage_5[14]), .I0( stage_4[14] ), .I1( stage_4[15] ), .I2( select[0] ) ); defparam mux_5_14.INIT = 8'hca; //'
    LUT3 mux_5_15 ( .O(stage_5[15]), .I0( stage_4[15] ), .I1( stage_4[16] ), .I2( select[0] ) ); defparam mux_5_15.INIT = 8'hca; //'
    LUT3 mux_5_16 ( .O(stage_5[16]), .I0( stage_4[16] ), .I1( stage_4[17] ), .I2( select[0] ) ); defparam mux_5_16.INIT = 8'hca; //'
    LUT3 mux_5_17 ( .O(stage_5[17]), .I0( stage_4[17] ), .I1( stage_4[18] ), .I2( select[0] ) ); defparam mux_5_17.INIT = 8'hca; //'
    LUT3 mux_5_18 ( .O(stage_5[18]), .I0( stage_4[18] ), .I1( stage_4[19] ), .I2( select[0] ) ); defparam mux_5_18.INIT = 8'hca; //'
    LUT3 mux_5_19 ( .O(stage_5[19]), .I0( stage_4[19] ), .I1( stage_4[20] ), .I2( select[0] ) ); defparam mux_5_19.INIT = 8'hca; //'
    LUT3 mux_5_20 ( .O(stage_5[20]), .I0( stage_4[20] ), .I1( stage_4[21] ), .I2( select[0] ) ); defparam mux_5_20.INIT = 8'hca; //'
    LUT3 mux_5_21 ( .O(stage_5[21]), .I0( stage_4[21] ), .I1( stage_4[22] ), .I2( select[0] ) ); defparam mux_5_21.INIT = 8'hca; //'
    LUT3 mux_5_22 ( .O(stage_5[22]), .I0( stage_4[22] ), .I1( stage_4[23] ), .I2( select[0] ) ); defparam mux_5_22.INIT = 8'hca; //'
    LUT3 mux_5_23 ( .O(stage_5[23]), .I0( stage_4[23] ), .I1( stage_4[24] ), .I2( select[0] ) ); defparam mux_5_23.INIT = 8'hca; //'
    LUT3 mux_5_24 ( .O(stage_5[24]), .I0( stage_4[24] ), .I1( stage_4[25] ), .I2( select[0] ) ); defparam mux_5_24.INIT = 8'hca; //'
    LUT3 mux_5_25 ( .O(stage_5[25]), .I0( stage_4[25] ), .I1( stage_4[26] ), .I2( select[0] ) ); defparam mux_5_25.INIT = 8'hca; //'
    LUT3 mux_5_26 ( .O(stage_5[26]), .I0( stage_4[26] ), .I1( stage_4[27] ), .I2( select[0] ) ); defparam mux_5_26.INIT = 8'hca; //'
    LUT3 mux_5_27 ( .O(stage_5[27]), .I0( stage_4[27] ), .I1( stage_4[28] ), .I2( select[0] ) ); defparam mux_5_27.INIT = 8'hca; //'
    LUT3 mux_5_28 ( .O(stage_5[28]), .I0( stage_4[28] ), .I1( stage_4[29] ), .I2( select[0] ) ); defparam mux_5_28.INIT = 8'hca; //'
    LUT3 mux_5_29 ( .O(stage_5[29]), .I0( stage_4[29] ), .I1( stage_4[30] ), .I2( select[0] ) ); defparam mux_5_29.INIT = 8'hca; //'
    LUT3 mux_5_30 ( .O(stage_5[30]), .I0( stage_4[30] ), .I1( stage_4[31] ), .I2( select[0] ) ); defparam mux_5_30.INIT = 8'hca; //'
    LUT3 mux_5_31 ( .O(stage_5[31]), .I0( stage_4[31] ), .I1( stage_4[ 0] ), .I2( select[0] ) ); defparam mux_5_31.INIT = 8'hca; //'

    assign out = stage_5;

endmodule
