/*a Includes
 */
include "gip.h"
include "gip_internal.h"

/*a Types
 */

/*a Module
 */
module gip_memory( clock gip_clock,
                   input bit gip_reset,

                   input t_gip_ins_r alu_mem_rd,
                   input bit mem_alu_busy,

                   output t_gip_ins_r mem_1_rd,
                   output t_gip_ins_r mem_2_rd,
                   input bit mem_read_data_valid
    )
"
    The GIP core memory stage is basically a simple pipeline; it is not responsible for delivering data, just tracking the external memory interface

    Basically it takes memory operation, and pushes them in to its pipe.

    It moves items down the pipeline, flowing them out when the external memory stage indicates the data is ready.
"

{

    /*b Clock and reset
     */
    default clock gip_clock;
    default reset gip_reset;

    /*b Pipeline
     */
    clocked t_gip_ins_r mem_1_rd = {type=gip_ins_r_type_none, r=0};
    clocked t_gip_ins_r mem_2_rd = {type=gip_ins_r_type_none, r=0};

    /*b Combinatorials
     */
    comb bit mem2_will_take_mem1 "This is asserted if mem2 is none, or if mem2 mem_read_data_valid is asserted";

    /*b Pipeline logic
     */
    pipeline "Pipeline the memory RDs":
        {
            mem2_will_take_mem1 = 0;
            if (mem_2_rd.type == gip_ins_r_type_none) // If the slot is empty, we will move up mem1
            {
                mem2_will_take_mem1 = 1;
            }
            if (mem_read_data_valid) // In this case we are returning data for the mem2 register
            {
                mem2_will_take_mem1 = 1;
            }
            
            if ( (alu_mem_rd.type != gip_ins_r_type_none) &&
                 !mem_alu_busy ) // If a read transaction is being taken by the memory then its register must be recorded
            {
                mem_1_rd <= alu_mem_rd;
            }
            else
            {
                if (mem2_will_take_mem1)
                {
                    mem_1_rd.type <= gip_ins_r_type_none;
                }
            }

            if (mem2_will_take_mem1)
            {
                mem_2_rd <= mem_1_rd;
            }
        }
}

