/*a Includes
 */
include "gip.h"

/*a Types
 */
/*t t_sram_data_op
 */
typedef enum [3]
{
    sram_data_op_word,
    sram_data_op_byte_0,
    sram_data_op_byte_1,
    sram_data_op_byte_2,
    sram_data_op_byte_3
} t_sram_data_op;

/*a Module
 */
module gip_data_ram( clock gip_clock,
                     input bit gip_reset,

                        input t_gip_mem_op alu_mem_op,
                        input t_gip_word alu_mem_address,
                        input t_gip_word alu_mem_write_data,
                        input bit[4] alu_mem_burst,

                        output bit mem_alu_busy,
                        output bit mem_read_data_valid,
                     output bit[32] mem_read_data,

                     output bit sram_not_in_use,
                     output bit sram_read_not_write,
                     output bit[4] sram_write_byte_enables,
                     output bit[32] sram_address,
                     output bit[32] sram_write_data,
                     input bit[32] sram_read_data

    )
"
    This data_ram model supports a simple model for the data memory for the GIP

    It can be shared with the instruction memory using the 'sram_not_in_use' output

    Basically operations are given to the data memory, which always takes them.
    The next cycle is the address cycle for the memory.
    The final cycle is the data cycle for the memory.

    This module is responsible for byte laning. It should have knowledge of accesses that are unaligned, also; but these are not supported here.
"

{

    /*b Clock and reset
     */
    default clock gip_clock;
    default reset gip_reset;

    /*b Outputs to the GIP core
     */
    clocked bit mem_alu_busy = 0;
    clocked bit mem_read_data_valid = 0;
    
    /*b SRAM interface
     */
    clocked bit sram_not_in_use = 0;
    clocked bit sram_read_not_write = 0;
    clocked bit[4] sram_write_byte_enables = 0;
    clocked bit[32] sram_address = 0;
    clocked bit[32] sram_write_data = 0;
    clocked t_sram_data_op sram_data_op = sram_data_op_word;
    clocked t_sram_data_op last_sram_data_op = sram_data_op_word;

    /*b SRAM interface code
     */
    sram_interface "SRAM interface":
        {
            sram_not_in_use <= 1;
            full_switch (alu_mem_op)
                {
                case gip_mem_op_none:
                {
                    sram_not_in_use <= 1;
                    sram_read_not_write <= 0;
                    sram_write_byte_enables <= 0;
                }
                case gip_mem_op_store_word:
                {
                    sram_not_in_use <= 0;
                    sram_read_not_write <= 0;
                    sram_write_byte_enables <= 15;
                    sram_write_data <= alu_mem_write_data;
                    sram_address <= alu_mem_address;
                }
                case gip_mem_op_store_byte:
                {
                    sram_not_in_use <= 0;
                    sram_read_not_write <= 0;
                    sram_write_byte_enables <= 0;
                    sram_write_byte_enables[alu_mem_address[2;0]] <= 1; // little endian
                    sram_write_data[8;0] <= alu_mem_write_data[8;0];
                    sram_write_data[8;8] <= alu_mem_write_data[8;0];
                    sram_write_data[8;16] <= alu_mem_write_data[8;0];
                    sram_write_data[8;24] <= alu_mem_write_data[8;0];
                    sram_address <= alu_mem_address;
                }
                case gip_mem_op_load_word:
                case gip_mem_op_load_byte:
                {
                    sram_not_in_use <= 0;
                    sram_read_not_write <= 1;
                    sram_write_byte_enables <= 0;
                    sram_address <= alu_mem_address;
                    sram_data_op <= sram_data_op_word;
                    if (alu_mem_op==gip_mem_op_load_byte)
                    {
                        full_switch (alu_mem_address[2;0])
                            {
                            case 0: {sram_data_op <= sram_data_op_byte_0; } // little endian
                            case 1: {sram_data_op <= sram_data_op_byte_1; } // little endian
                            case 2: {sram_data_op <= sram_data_op_byte_2; } // little endian
                            case 3: {sram_data_op <= sram_data_op_byte_3; } // little endian
                            }
                    }
                }
                }
        }

    /*b GIP interface
     */
    gip_interface "GIP interface code":
        {
            mem_read_data = 0;
            full_switch (last_sram_data_op)
                {
                case sram_data_op_word:
                {
                    mem_read_data = sram_read_data;
                }
                case sram_data_op_byte_0:
                {
                    mem_read_data[8;0] = sram_read_data[8;0];
                }
                case sram_data_op_byte_1:
                {
                    mem_read_data[8;0] = sram_read_data[8;8];
                }
                case sram_data_op_byte_2:
                {
                    mem_read_data[8;0] = sram_read_data[8;16];
                }
                case sram_data_op_byte_3:
                {
                    mem_read_data[8;0] = sram_read_data[8;24];
                }
                }
            last_sram_data_op <= sram_data_op;
            mem_read_data_valid <= sram_read_not_write;
            mem_alu_busy <= 0;
        }
}
