/*a Copyright Gavin J Stark, 2004
 */

/*a Includes
 */
include "io_uart.h"
include "apb_target_uart.h"
include "apb_target_ext_bus_master.h"
include "apb_target_gpio.h"
include "apb_target_timer.h"

/*a Types
 */
/*t t_global_apb_state
 */
typedef fsm
{
    global_apb_state_idle         "APB idle";
    global_apb_state_write_select "APB writing, select asserted, no enable";
    global_apb_state_write_enable "APB writing, select and enable asserted";
    global_apb_state_read_select  "APB reading, select asserted, no enable";
    global_apb_state_read_enable  "APB reading, select and enable asserted, data should be valid (unless wait asserted)";
    global_apb_state_recover      "APB done reading/writing; read data valid to internal APB, write just waiting for enable to go away";
} t_global_apb_state;

/*a Modules
 */
module apb_devices( clock int_clock,
                    input bit int_reset,

                    input bit apb_pselect,
                    input bit apb_penable,
                    input bit apb_prnw,
                    input bit[6] apb_paddr,
                    input bit[32] apb_pwdata,
                    output bit[32] apb_prdata,
                    output bit apb_pwait,

                    output bit global_apb_pselect,
                    output bit global_apb_penable,
                    output bit global_apb_prnw,
                    output bit[5] global_apb_paddr,
                    output bit[32] global_apb_pwdata,
                    input bit[32] global_apb_prdata,
                    input bit global_apb_pwait,

                    output bit txd,
                    input bit rxd,
                    output bit[4]ext_bus_ce,
                    output bit ext_bus_oe,
                    output bit ext_bus_we,
                    output bit[24]ext_bus_address,
                    output bit ext_bus_write_data_enable,
                    output bit[32]ext_bus_write_data,
                    input bit[32]ext_bus_read_data,

                    input bit[4]gpio_input,
                    output bit[16]gpio_output,
                    output bit[16]gpio_output_enable,
                    output bit gpio_input_event,

                    output bit[3] timer_equalled
    )
{
    default clock int_clock;
    default reset int_reset;

    net bit[4]ext_bus_ce;
    net bit ext_bus_oe;
    net bit ext_bus_we;
    net bit[24]ext_bus_address;
    net bit ext_bus_write_data_enable;
    net bit[32]ext_bus_write_data;

    comb bit tx_baud_enable "Baud enable for transmit, 16 x bit time";
    net bit txd "Transmit data out";
//    net bit txd_fc "Transmit flow control; assert to pause transmit";

    comb bit rx_baud_enable "Baud enable for receive, 16 x bit time";
    net bit rxd_fc "Receive flow control; asserted to pause transmit";

    net bit cmd_fifo_empty;
    net bit[32] cmd_fifo_data;
    net bit cmd_fifo_toggle;

    net bit status_fifo_full;
    net bit status_fifo_toggle;
    net bit[32] status_fifo_data;

    net bit[32] apb_prdata_uart;
    net bit[32] apb_prdata_ext_bus;
    net bit[32] apb_prdata_gpio;
    net bit[32] apb_prdata_timer;
    clocked bit[32] apb_prdata_global = 0;
    net bit apb_pwait_ext_bus;
    net bit apb_pwait_timer;
    comb bit apb_pwait_global;
    clocked t_global_apb_state global_apb_state = global_apb_state_idle;
    clocked bit[32] global_apb_pwdata = 0;
    clocked bit[5] global_apb_paddr = 0;

    comb bit[2] cfg_uart_speed;
    comb bit[16] cfg_baud_divider;
    clocked bit[16] baud_counter=0;
    clocked bit[6] baud_divider = 0;

    net bit[16]gpio_output;
    net bit[16]gpio_output_enable;
    net bit gpio_input_event;
    net bit[3] timer_equalled;

    /*b Clock divider
     */
    divider "Clock divider for LED":
        {
            cfg_uart_speed = 0;
            full_switch( cfg_uart_speed )
                {
                case 0: // 260=>9600 - actually 1200 for 5MHz; for 125/12 we need 60
                {
                    cfg_baud_divider = 260;
                    cfg_baud_divider = 68;
                }
                case 1: // 130=>19200 - actually 2400 for 5MHz and for 125/12 we need 241
                {
                    cfg_baud_divider = 130;
                    cfg_baud_divider = 271;
                }
                case 2: // 38400 - NOW 10Hz for 5MHz
                {
                    cfg_baud_divider = 65;
                    cfg_baud_divider = 16h7a21; // 31250 = 5,000,000/160
                    cfg_baud_divider = 34;
                }
                case 3: // none - i.e. divide by 8
                {
                    cfg_baud_divider = 8;
                }
                }
            baud_counter <= baud_counter+1;
            if (baud_counter+1 == cfg_baud_divider)
            {
                baud_counter <= 0;
            }
            rx_baud_enable = (baud_counter==0);
            tx_baud_enable = rx_baud_enable;
            if (rx_baud_enable)
            {
                baud_divider <= baud_divider+1;
            }
        }

    /*b APB instances
     */
    apb_instances "APB Instances":
        {
            apb_target_uart uart_apb( apb_clock <- int_clock,
                                      int_reset <= int_reset,

                                      apb_pselect <= apb_pselect && (apb_paddr[3;3]==0),
                                      apb_penable <= apb_penable,
                                      apb_paddr <= apb_paddr[3;0],
                                      apb_prnw <= apb_prnw,
                                      apb_pwdata <= apb_pwdata,
                                      apb_prdata => apb_prdata_uart,
                                      
                                      cmd_fifo_empty => cmd_fifo_empty,
                                      cmd_fifo_data => cmd_fifo_data,
                                      cmd_fifo_toggle <= cmd_fifo_toggle,

                                      status_fifo_full => status_fifo_full,
                                      status_fifo_data <= status_fifo_data,
                                      status_fifo_toggle <= status_fifo_toggle );

            apb_target_ext_bus_master ext_bus_apb( apb_clock <- int_clock,
                                                   int_reset <= int_reset,

                                                   apb_pselect <= apb_pselect && (apb_paddr[3;3]==1),
                                                   apb_penable <= apb_penable,
                                                   apb_paddr <= apb_paddr[3;0],
                                                   apb_prnw <= apb_prnw,
                                                   apb_pwdata <= apb_pwdata,
                                                   apb_prdata => apb_prdata_ext_bus,
                                                   apb_pwait => apb_pwait_ext_bus,

                                                   ext_bus_ce => ext_bus_ce,
                                                   ext_bus_oe => ext_bus_oe,
                                                   ext_bus_we => ext_bus_we,
                                                   ext_bus_address => ext_bus_address,
                                                   ext_bus_write_data_enable => ext_bus_write_data_enable,
                                                   ext_bus_write_data => ext_bus_write_data,
                                                   ext_bus_read_data <= ext_bus_read_data );

            apb_target_gpio gpio_apb( apb_clock <- int_clock,
                                      int_reset <= int_reset,

                                      apb_pselect <= apb_pselect && (apb_paddr[3;3]==2),
                                      apb_penable <= apb_penable,
                                      apb_paddr <= apb_paddr[3;0],
                                      apb_prnw <= apb_prnw,
                                      apb_pwdata <= apb_pwdata,
                                      apb_prdata => apb_prdata_gpio,

                                      gpio_output => gpio_output,
                                      gpio_output_enable => gpio_output_enable,
                                      gpio_input <= gpio_input,
                                      gpio_input_event => gpio_input_event );

            apb_target_timer timer_apb( apb_clock <- int_clock,
                                        int_reset <= int_reset,

                                        apb_pselect <= apb_pselect && (apb_paddr[3;3]==3),
                                        apb_penable <= apb_penable,
                                        apb_paddr <= apb_paddr[3;0],
                                        apb_prnw <= apb_prnw,
                                        apb_pwdata <= apb_pwdata,
                                        apb_prdata => apb_prdata_timer,
                                        apb_pwait => apb_pwait_timer,

                                        timer_equalled => timer_equalled );

            full_switch (apb_paddr[3;3])
                {
                case 0:  {apb_prdata = apb_prdata_uart;    apb_pwait = 0;}
                case 1:  {apb_prdata = apb_prdata_ext_bus; apb_pwait = apb_pwait_ext_bus;}
                case 2:  {apb_prdata = apb_prdata_gpio;    apb_pwait = 0;}
                case 3:  {apb_prdata = apb_prdata_timer;   apb_pwait = apb_pwait_timer;}
                default: {apb_prdata = apb_prdata_global;  apb_pwait = apb_pwait_global;}
                }
        }

    /*b Global APB FSM
     */
    global_apb_state_machine "FSM and decode for global APB":
        {
            global_apb_paddr <= apb_paddr[5;0];
            global_apb_pselect = 0;
            global_apb_penable = 0;
            global_apb_prnw = 0;
            apb_pwait_global = 0;
            full_switch (global_apb_state)
                {
                case global_apb_state_idle:
                {
                    global_apb_pselect = 0;
                    global_apb_penable = 0;
                    global_apb_prnw = 0;
                    apb_pwait_global = 0;
                    if (apb_pselect && apb_paddr[5]) // if global
                    {
                        if (apb_prnw)
                        {
                            global_apb_state <= global_apb_state_read_select;
                        }
                        else
                        {
                            global_apb_state <= global_apb_state_write_select;
                            global_apb_pwdata <= apb_pwdata;
                        }
                    }
                }
                case global_apb_state_read_select: // internal apb will be presenting enable, we need to hold that until we have data in our buffer
                {
                    global_apb_pselect = 1;
                    global_apb_penable = 0;
                    global_apb_prnw = 1;
                    apb_pwait_global = 1;
                    if (!global_apb_pwait)
                    {
                        global_apb_state <= global_apb_state_read_enable;
                    }
                }
                case global_apb_state_read_enable: // internal apb will be presenting enable, we need to hold that until we have data in our buffer
                {
                    global_apb_pselect = 1;
                    global_apb_penable = 1;
                    global_apb_prnw = 1;
                    apb_pwait_global = 1;
                    if (!global_apb_pwait)
                    {
                        global_apb_state <= global_apb_state_recover;
                        apb_prdata_global <= global_apb_prdata;
                    }
                }
                case global_apb_state_write_select: // internal apb will be presenting enable, we need to hold APB and present select to global APB (we cannot let internal APB run as it may do another transaction!)
                {
                    global_apb_pselect = 1;
                    global_apb_penable = 0;
                    global_apb_prnw = 0;
                    apb_pwait_global = 1;
                    if (!global_apb_pwait)
                    {
                        global_apb_state <= global_apb_state_write_enable;
                    }
                }
                case global_apb_state_write_enable: // internal apb will be presenting enable, we need to hold APB and present enable to global APB (we cannot let internal APB run as it may do another transaction!)
                {
                    global_apb_pselect = 1;
                    global_apb_penable = 1;
                    global_apb_prnw = 0;
                    apb_pwait_global = 1;
                    if (!global_apb_pwait)
                    {
                        global_apb_state <= global_apb_state_recover; // ensure that we enter idle with the current transaction just complete
                    }
                }
                case global_apb_state_recover: // internal apb will be presenting enable, and for reads we have the read data to present, for writes we just need to wait
                {
                    global_apb_pselect = 0;
                    global_apb_penable = 0;
                    global_apb_prnw = 0;
                    apb_pwait_global = 0;
                    global_apb_state <= global_apb_state_idle;
                }
                }
        }

    /*b Extra components for APB-based IO UART
     */
    uart_comps "Extra components for APB-based IO UART":
        {
            io_uart uart_io( int_clock <- int_clock,
                          int_reset <= int_reset,
                          tx_baud_enable <= tx_baud_enable,
                          txd => txd,
                          txd_fc <= 0,
                          rx_baud_enable <= rx_baud_enable,
                          rxd <= rxd,
                          rxd_fc => rxd_fc,

                          cmd_fifo_empty <= cmd_fifo_empty,
                          cmd_fifo_data <= cmd_fifo_data,
                          cmd_fifo_toggle => cmd_fifo_toggle,

                          status_fifo_full <= status_fifo_full,
                          status_fifo_data => status_fifo_data,
                          status_fifo_toggle => status_fifo_toggle );

        }

}

