/*a Copyright Gavin J Stark, 2004
 */

/*a To do
Ensure status is writing time and data to successive locations
 */

/*a Includes
 */
include "io_cmd.h"
include "io.h"
include "postbus.h"

include "io_ethernet_rx.h"
include "io_ethernet_tx.h"
include "io_sync_serial.h"
include "io_uart.h"
include "io_baud_rate_generator.h"

include "io_sync_request.h"
include "io_ingress_fifos.h"
include "io_egress_fifos.h"
include "io_egress_control.h"
include "io_ingress_control.h"
include "io_postbus.h"
include "memories.h"

/*a Constants
 */

/*a Types
 */
/*t t_postbus_src_read_data_source
 */
typedef enum [2]
{
    postbus_src_read_data_source_ingress_fifo_status,
    postbus_src_read_data_source_ingress_sram,
    postbus_src_read_data_source_egress_fifo_status,
    postbus_src_read_data_source_egress_sram,
} t_postbus_src_read_data_source;

/*t t_io_port_config
 */
typedef struct
{
    bit in_reset; // if 1, inputs are ignored from the port - also this signal goes to the port as a reset signal
    bit[2] fifo; // fifos to use for this port
    bit little_endian; // if 1 then network data FIFO data is byte swapped, as it network interfaces are assumed to be byte-wise and use/fill data words in a big endian manner
    bit[2] config; // config for the interface itself
} t_io_port_config;

/*a io_block module
 */
module io_block( clock int_clock,
                 input bit int_reset,

                 input t_postbus_type postbus_tgt_type "Postbus target bus type",
                 input t_postbus_data postbus_tgt_data "Postbus target bus data",
                 output t_postbus_ack postbus_tgt_ack  "Postbus target bus ack",

                 output t_postbus_type postbus_src_type  "Postbus source bus type",
                 output t_postbus_data postbus_src_data  "Postbus source bus data",
                 input t_postbus_ack postbus_src_ack     "Postbus source bus ack",

                 output bit    io_slot_cfg_write "asserted if cfg_data should be written to cfg_slot",
                 output bit[8] io_slot_cfg_data  "data for setting a slot configuration",
                 output bit[2] io_slot_cfg_slot  "number of slot cfg data is destined for",

                 input bit[4]    io_slot_egr_cmd_ready  "bus of command emptys from all slots - they are filled asynchronously to requests",
                 input bit       io_slot_egr_data_req    "OR of data requests, masked by pending acknowledgements",
                 input t_io_tx_data_fifo_cmd   io_slot_egr_data_cmd    "data command from lowest number slot with an unmasked request",
                 input bit[2]    io_slot_egr_data_slot   "slot the data command is coming from",
                 output bit      io_slot_egr_data_ack "asserted to acknowledge the current data request",
                 output bit[32]  io_slot_egr_data "contains data for writes to the slots, registered here, valid 3 cycles after acknowledged request (acked req in cycle 0, sram req in cycle 1, sram data stored end cycle 2, this valid in cycle 3",
                 output bit[2]   io_slot_egr_slot "indicates which slot the egress data is for, registered here; ",
                 output bit      io_slot_egr_cmd_write  "asserted if the data on the bus in this cycle is for the command side interface - if so, it will drive the not empty signal to the slot client",
                 output bit      io_slot_egr_data_write "asserted if the data on the bus in this cycle is for the data side interface",

                 input bit[32]  io_slot_ingr_data       "muxed in slot head from clients, ANDed with a select from io_slot_ing_number",
                 input bit      io_slot_ingr_status_req "OR of status requests, masked by pending acknowledgements",
                 input bit      io_slot_ingr_data_req    "OR of rx data requests, masked by pending acknowledgements, clear if status_req is asserted",
                 input bit[2]   io_slot_ingr_slot       "indicates which slot the status or rx data request is from",
                 output bit     io_slot_ingr_ack        "acknowledge, valid in same clock as status_req and data_req",
                 output bit[4]  io_slot_ingr_data_full  "for use by I/O",

                 input bit[3] analyzer_mux_control "Logic analyzer multiplex control, registered internally",
                 output bit[32] analyzer_signals   "Logic analyzer output signals, registered internally"
    )

    /*b Documentation
     */
"
This basically consists of a postbus interface to two main I/O subsections, ingress and egress, and the interfaces attached to the ingress and egress

Ingress and egress each have a 2kB by 32 bit RAM that implements a command/status set of 4 FIFOs and a set of 4 data FIFOs.

Each I/O interface then attaches to one of the four slots; the I/O interface should have a command interface for 32-bit commands to the interface, a status interface for 32-bit status indications, and they may also use a transmit data FIFO and/or a received data FIFO.

The I/O interfaces receive 'not empty' indications for commands and transmit data, but these have different semantics.
The command 'not empty' means that the command data is sitting on the bus in to the I/O interface, and acknowledging the command results in it changing.
The tx data 'not empty' means that transmit data can be fetched from the data FIFO; a command must then be issued to make the data appear, with a request.

The status and rx data FIFOs operate by presenting data with a request.

The synchronization for these interfaces is novel. Each request is presented by toggling a signal; this toggle is synchronized to the internal clock domain, which handles the requests from the active I/O interfaces.
The internal clock domain handles the requests in priority order (interface 0 through 3), intermixing with single words from the postbus side, so a request from interface 0 for transmit data takes up to 3 internal cycles for synchronization, one for request preparation, one for presentation to SRAM, one to perform an SRAM access, one to transfer the data to the slot head, then another to present the data; this is a total of 8 internal cycles plus data routing time. The requests from the I/O interface, therefore, must be placed at least 8 internal cycles apart, which would mean that for 8-bit wide I/O interfaces they must run at slower than internal clock/8*4.

The same restrictions apply to the status and receive data, with the caveat that receive status actually requires two internal clocks to write a time and a status indication word, so it requires 8 internal cycles of holdoff between the request and the status data from the interface changing or the status request toggling again.

For interfaces with lower priority the constraints of the higher priority interface should feed in to their calculations. Usually this is irrelevant, as the rate of requests from an interface will be less than one per 8 cycles, which should allow space for almost peak rates for each interface; but the actual latency should be increased by 4 internal cycles per interface, for safe operation.

The command interface consists of:
  dirn      signal    size   clock   description
to I/O      empty       1     int    brought low to indicate the command data bus has valid data - should be synchronized to i/o clock domain
from I/O    toggle      1     i/o    toggled to indicate acknowledgement of a valid command on the command data pins; after this toggles, the command data should be deemed invalid; the empty signal will assert after at most 4 internal clock ticks
to I/O      data       32     int    always qualify with a synchronized empty signal so the data need not be synchronized

The tx data interface consists of:
  dirn      signal    size   clock   description
from I/O    cmd       cmd     i/o    indicates read, read and commit, commit, or revert
from I/O    toggle      1     i/o    toggled to indicate request for the corresponding command to occur
to I/O      data       32     int    presents data read in response to a read command, at 8+ internal clocks after the command

The rx data interface consists of:
  dirn      signal    size   clock   description
to I/O      full        1     int    indicates the receive data FIFO is full - asserted when a write takes place filling the FIFO. May be used (synchronized) to effect operation of the I/O.
from I/O    toggle      1     i/o    toggled to indicate request for data to be written to the FIFO
from I/O    data       32     i/o    contains data to be written to the receive data FIFO; must be stable for 8+ internal clocks after the toggle

The rx status interface consists of:
  dirn      signal    size   clock   description
to I/O      full        1     int    indicates the receive status FIFO is full - asserted when a write takes place filling the FIFO. May be used (synchronized) to effect operation of the I/O.
from I/O    toggle      1     i/o    toggled to indicate request for status to be written to the FIFO
from I/O    data       32     i/o    contains data to be written to the receive status FIFO; must be stable for 8+ internal clocks after the toggle


A standard module (io_sync_request) is used to synchronize the toggle signals to generate internal requests, which are acknowledged also off the internal clock domain.

We have in each module:
2 ethernet (tx plus rx)
2 general purpose (flexible I/O)
1 async serial
1 sync serial (MDIO/SPI)
1 usb

Slot 0 is always ethernet A
Slot 1 is either ethernet B or a general purpose data in/out A
Slot 2 is either sync serial of general purpose data in/out B
Slot 3 is either async serial or USB

Each interface slot requires its own io_sync_request modules for each of the toggles.
For data to the I/O, each slot has a register which stores the command or data, and it drives all the interfaces which may be attached to that slot; the main block drives the data out from a register with controls indicating which slot it is for.
For data (rx status and rx data) and cmd (tx data) from the I/O, these are ORed together at the slot head
Each slot also has 8 control signal associated with it, which may be used to reset the various interfaces attached to the slot, and indicate which client of the slot is selected.

So this level has...


to I/O     io_slot_cfg_data (contains data for setting a slot configuration)
to I/O     io_slot_cfg_slot (number of slot cfg data is destined for)
to I/O     io_slot_cfg_write (asserted if cfg_data should be written

from I/O   io_slot_egr_cmd_empty (bus of command emptys from all slots - they are filled asynchronously to requests)
from I/O   io_slot_egr_data_req (OR of data requests, masked by pending acknowledgements)
from I/O   io_slot_egr_data_cmd (data command from lowest number slot with an unmasked request)
from I/O   io_slot_egr_data_slot (slot the data command is coming from)

to I/O     io_slot_egr_data (contains data for writes to the slots, registered here, valid 3 cycles after acknowledged request (acked req in cycle 0, sram req in cycle 1, sram data stored end cycle 2, this valid in cycle 3)
to I/O     io_slot_egr_slot (indicates which slot the egress data is for, registered here; )
to I/O     io_slot_egr_cmd_not_data (asserted if the data on the bus in this cycle is for the command side interface - if so, it will drive the not empty signal to the slot client)

from I/O   io_slot_ingr_data (muxed in slot head from clients, ANDed with a select from io_slot_ing_number)
from I/O   io_slot_ingr_status_req (OR of status requests, masked by pending acknowledgements)
from I/O   io_slot_ingr_rxd_req    (OR of rx data requests, masked by pending acknowledgements, clear if status_req is asserted)
from I/O   io_slot_ingr_slot       (indicates which slot the status or rx data request is from)
to I/O     io_slot_ingr_ack        (acknowledge, valid in same clock as status_req and rxd_req)
to I/O     io_slot_ingr_data_full  (for use by the I/O)
"
{

    /*b -------------------- Registers, nets and combinatorials
     */

    /*b Default clock and reset - internal clock domain
     */
    default clock int_clock;
    default reset int_reset;

    /*b Logic analyzer control
     */
    clocked bit[3] analyzer_mux_control_reg = 0 "Register the analyzer mux control to reduce any timing issues on this bus system";
    clocked bit[32] analyzer_signals = 0 "Registered logic analyzer output signals, registered internally to reduce any timing issues on the bus system";

    /*b I/O Slot registers
     */
    clocked bit io_slot_cfg_write = 0;
    clocked bit[2] io_slot_cfg_slot = 0;
    clocked bit[8] io_slot_cfg_data = 0;

//    clocked bit io_slot_egr_data_ack "asserted to acknowledge the current data request",
    clocked bit[32]  io_slot_egr_data = 0;
    clocked bit[2]   io_slot_egr_slot = 0;
    clocked bit      io_slot_egr_cmd_write  = 0;
    clocked bit      io_slot_egr_data_write = 0;

    clocked bit rx_data_req = 0;
    clocked bit status_req = 0;
    clocked bit io_slot_ingr_ack = 0;
    net bit status_rx_data_will_be_acked;
    clocked bit[2] status_rx_data_fifo = 0;
    clocked bit[32] status_rx_data_fifo_data = 0;

    clocked bit[4] cmd_available_bus = 0;
    net bit        cmd_valid "Asserted if the SRAM has a command for a slot";
    net bit[2]     cmd_valid_number "If cmd_valid is asserted, then it indicates which slot the command is for";

    clocked bit    tx_data_req = 0     "Asserted if we are requesting data for one of the slots";
    net bit tx_data_ack;
    clocked bit[2] tx_data_req_num = 0 "Number of the slot we are requesting data for";
    clocked t_io_tx_data_fifo_cmd tx_data_cmd = io_tx_data_fifo_cmd_read_fifo "Command to do if request asserted";

    clocked bit[4] last_io_slot_egr_cmd_ready = 0;

    clocked bit tx_data_read_being_presented=0;
    clocked bit[2] tx_data_slot_being_presented=0;
    clocked bit tx_data_reading = 0;
    clocked bit[2] tx_data_slot_reading = 0;

    /*b Ingress arbiter and controller wiring
     */
    net bit ingress_postbus_req;
    net bit ingress_postbus_ack;

    net t_io_sram_data_op ingress_sram_data_op;
    net bit ingress_sram_data_reg_hold;
    net t_io_sram_address_op ingress_sram_address_op;

    net t_io_fifo_op ingress_fifo_op;
    net bit ingress_fifo_op_to_status;
    net bit[2] ingress_fifo_to_access;
    net bit ingress_fifo_address_from_read_ptr;
    net t_io_fifo_event_type ingress_fifo_event_type;
    net bit[io_sram_log_size] ingress_fifo_address;
    net bit[32] ingress_fifo_cfg_status;
    net bit ingress_event_from_status;
    net bit[2] ingress_event_fifo;
    net t_io_fifo_event ingress_event_empty;
    net t_io_fifo_event ingress_event_watermark;

    clocked bit[32] ingress_data_reg = 0;

    /*b Egress arbiter and controller wiring
     */
    net bit egress_postbus_req;
    net bit egress_postbus_ack;

    net t_io_sram_data_op egress_sram_data_op;
    net t_io_sram_data_reg_op egress_sram_data_reg_op;
    net t_io_sram_address_op egress_sram_address_op;

    net t_io_fifo_op egress_fifo_op;
    net bit egress_fifo_op_to_cmd;
    net bit[2] egress_fifo_to_access;
    net bit egress_fifo_address_from_read_ptr;
    net t_io_fifo_event_type egress_fifo_event_type;
    net bit[io_sram_log_size] egress_fifo_address;
    net bit[32] egress_fifo_cfg_status;
    net bit egress_event_from_cmd;
    net bit[2] egress_event_fifo;
    net t_io_fifo_event egress_event_empty;
    net t_io_fifo_event egress_event_watermark;

    clocked bit[32] egress_data_reg = 0;

    /*b Postbus registers
     */
    net t_postbus_ack postbus_tgt_ack;

    net t_postbus_type postbus_src_type;
    net t_postbus_data postbus_src_data;
    comb bit[32] postbus_src_read_data;

    net bit[32] postbus_write_data;
    net bit[5] postbus_write_address;
    net bit postbus_configuration_write;

    net t_io_fifo_op         egress_postbus_fifo_op;
    net bit                  egress_postbus_fifo_op_to_cmd_status;
    net bit[2]               egress_postbus_fifo_to_access;
    net t_io_fifo_event_type egress_postbus_fifo_event_type;
    net bit                  egress_postbus_fifo_address_from_read_ptr;
    net t_io_sram_address_op egress_postbus_sram_address_op;
    net t_io_sram_data_op    egress_postbus_sram_data_op;

    net t_io_fifo_op         ingress_postbus_fifo_op;
    net bit                  ingress_postbus_fifo_op_to_cmd_status;
    net bit[2]               ingress_postbus_fifo_to_access;
    net t_io_fifo_event_type ingress_postbus_fifo_event_type;
    net bit                  ingress_postbus_fifo_address_from_read_ptr;
    net t_io_sram_address_op ingress_postbus_sram_address_op;
    net t_io_sram_data_op    ingress_postbus_sram_data_op;

    clocked t_postbus_src_read_data_source postbus_src_read_data_source = postbus_src_read_data_source_egress_sram;
    clocked t_postbus_src_read_data_source next_postbus_src_read_data_source = postbus_src_read_data_source_egress_sram;
    clocked bit[32] sram_read_data_fifo_status = 0;

    /*b Status registers
     */
    clocked bit[32] status_timer = 0;

    /*b Ingress SRAM control signals
     */
    comb bit ingress_sram_write;
    comb bit ingress_sram_read;
    comb bit[io_sram_log_size] ingress_sram_address;
    comb bit[32] ingress_sram_write_data;
    net bit[32] ingress_sram_read_data;

    /*b Egress SRAM control signals
     */
    comb bit egress_sram_write;
    comb bit egress_sram_read;
    comb bit[io_sram_log_size] egress_sram_address;
    comb bit[32] egress_sram_write_data;
    net bit[32] egress_sram_read_data;

    /*b Fifo wiring
     */
    net bit[4] cmd_fifo_empty       "Per-cmd FIFO, asserted if more than zero entries are present";
    net bit[4] cmd_fifo_full        "Per-cmd FIFO, asserted if read_ptr==write_ptr and not empty";
    net bit[4] cmd_fifo_overflowed  "Per-cmd FIFO, asserted if FIFO has overflowed since last reset or configuration write";
    net bit[4] cmd_fifo_underflowed "Per-cmd FIFO, asserted if FIFO has underflowed since last reset or configuration write";

    net bit[4] status_fifo_empty       "Per-status FIFO, asserted if more than zero entries are present";
    net bit[4] status_fifo_full        "Per-status FIFO, asserted if read_ptr==write_ptr and not empty";
    net bit[4] status_fifo_overflowed  "Per-status FIFO, asserted if FIFO has overflowed since last reset or configuration write";
    net bit[4] status_fifo_underflowed "Per-status FIFO, asserted if FIFO has underflowed since last reset or configuration write";

    net bit[4] tx_data_fifo_empty       "Per-tx_data FIFO, asserted if more than zero entries are present";
    net bit[4] tx_data_fifo_watermark   "Per-tx_data FIFO, asserted if more than watermak entries are present in the FIFO";
    net bit[4] tx_data_fifo_full        "Per-tx_data FIFO, asserted if read_ptr==write_ptr and not empty";
    net bit[4] tx_data_fifo_overflowed  "Per-tx_data FIFO, asserted if FIFO has overflowed since last reset or configuration write";
    net bit[4] tx_data_fifo_underflowed "Per-tx_data FIFO, asserted if FIFO has underflowed since last reset or configuration write";

    net bit[4] rx_data_fifo_empty       "Per-rx_data FIFO, asserted if more than zero entries are present";
    net bit[4] rx_data_fifo_watermark   "Per-rx_data FIFO, asserted if more than watermak entries are present in the FIFO";
    net bit[4] rx_data_fifo_full        "Per-rx_data FIFO, asserted if read_ptr==write_ptr and not empty";
    net bit[4] rx_data_fifo_overflowed  "Per-rx_data FIFO, asserted if FIFO has overflowed since last reset or configuration write";
    net bit[4] rx_data_fifo_underflowed "Per-rx_data FIFO, asserted if FIFO has underflowed since last reset or configuration write";

    comb bit[io_sram_log_size] cfg_base_address;
    comb bit[io_sram_log_size] cfg_size_m_one;
    comb bit[io_sram_log_size] cfg_watermark;

    /*b Baud rate generator wiring
     */
    comb bit brg0_counter_enable "Assert to run BRG0";
    comb bit brg0_counter_reset "Assert to reset BRG0 counter, to sync multiple BRGs";
    net bit brg0_baud_enable "Output of BRG0";
    comb bit brg0_set_config "Assert to write config data to BRG0";

    comb bit brg1_counter_enable "Assert to run BRG1";
    comb bit brg1_counter_reset "Assert to reset BRG1 counter, to sync multiple BRGs";
    net bit brg1_baud_enable "Output of BRG1";
    comb bit brg1_set_config "Assert to write config data to BRG1";

    comb bit[io_baud_rate_divider_size] cfg_baud_addition_value;
    comb bit[io_baud_rate_divider_size] cfg_baud_subtraction_value;

    /*b -------------------- Logic
     */

    /*b Analyzer signals
     */
    analyzer_signal_setting "Analyzer signals":
        {
            analyzer_mux_control_reg <= analyzer_mux_control;
            analyzer_signals <= 0;
            part_switch (analyzer_mux_control_reg)
                {
                case 0: // egress sram signals
                {
                    analyzer_signals[0] <= egress_sram_write;
                    analyzer_signals[1] <= egress_sram_read;
                    analyzer_signals[2] <= egress_fifo_op_to_cmd;
                    analyzer_signals[2;3] <= egress_fifo_to_access;
                    analyzer_signals[3;5] <= egress_fifo_op;
                    analyzer_signals[8] <= egress_fifo_address_from_read_ptr;
                    analyzer_signals[2;9] <= egress_fifo_event_type;
                    analyzer_signals[11] <= egress_event_from_cmd;
                    analyzer_signals[2;12] <= egress_event_fifo;
                    analyzer_signals[14] <= egress_postbus_req;
                    analyzer_signals[15] <= egress_postbus_ack;
                    analyzer_signals[16] <= tx_data_req;
                    analyzer_signals[17] <= cmd_valid;
                    analyzer_signals[io_sram_log_size;18] <= egress_sram_address;
                }
                case 1: // ingress sram signals
                {
                    analyzer_signals[0] <= ingress_sram_write;
                    analyzer_signals[1] <= ingress_sram_read;
                    analyzer_signals[2] <= ingress_fifo_op_to_status;
                    analyzer_signals[2;3] <= ingress_fifo_to_access;
                    analyzer_signals[3;5] <= ingress_fifo_op;
                    analyzer_signals[8] <= ingress_fifo_address_from_read_ptr;
                    analyzer_signals[2;9] <= ingress_fifo_event_type;
                    analyzer_signals[11] <= ingress_event_from_status;
                    analyzer_signals[2;12] <= ingress_event_fifo;
                    analyzer_signals[14] <= ingress_postbus_req;
                    analyzer_signals[15] <= ingress_postbus_ack;
                    analyzer_signals[16] <= rx_data_req;
                    analyzer_signals[17] <= status_req;
                    analyzer_signals[io_sram_log_size;18] <= ingress_sram_address;
                }
                }
        }

    /*b IO status/rx data slot interface
     */
    io_status_rx_data_slot_interface "IO status and receive data slot interface":
        {
            // this interface works as follows:
            //       0              1             2                    3                   4             5
            // sreqin,ack   sreq,sreqin,ack  sreq,!ack,wrtime    sreq,ack,wrdata       !ack,wrtime      ack,wrdata
            //              srdfd status     dreg st, srdfd st2  dreg st, srdfd st2      dreg st2        dreg st2
            //
            //       0              1             2                    3                   4   
            // dreqin,ack   dreq,dreqin,ack  dreq,ack,wrdata   dreq,ack,wrdata       ack,wrdata
            //              srdfd data       dreg d, srdfd d2  dreg d2, srdfd d3      dreg d3
            if (io_slot_ingr_ack)
            {
                status_req <= io_slot_ingr_status_req;
                rx_data_req <= io_slot_ingr_data_req;
                status_rx_data_fifo <= io_slot_ingr_slot;
                status_rx_data_fifo_data <= io_slot_ingr_data;
            }
            io_slot_ingr_ack <= status_rx_data_will_be_acked;

            io_slot_ingr_data_full = rx_data_fifo_full;

        }

    /*b Status and RxData FIFO ptrs and their arbiter
     */
    status_fifos_and_arbiter "Status, Rx data fifos, and arbiter":
        {
            io_ingress_control ingress_control( int_clock <- int_clock,
                                                int_reset <= int_reset,
                                                status_req <= status_req,
                                                rx_data_req <= rx_data_req,
                                                status_rx_data_fifo <= status_rx_data_fifo,
                                                status_rx_data_will_be_acked => status_rx_data_will_be_acked,

                                                postbus_req <= ingress_postbus_req,
                                                postbus_ack => ingress_postbus_ack,

                                                postbus_fifo_op <= ingress_postbus_fifo_op,
                                                postbus_fifo_address_from_read_ptr <= ingress_postbus_fifo_address_from_read_ptr,
                                                postbus_fifo_op_to_status <= ingress_postbus_fifo_op_to_cmd_status,
                                                postbus_fifo_event_type <= ingress_postbus_fifo_event_type,
                                                postbus_fifo_to_access <= ingress_postbus_fifo_to_access,

                                                postbus_sram_data_op <= ingress_postbus_sram_data_op,
                                                postbus_sram_address_op <= ingress_postbus_sram_address_op,

                                                ingress_fifo_op => ingress_fifo_op,
                                                ingress_fifo_op_to_status => ingress_fifo_op_to_status,
                                                ingress_fifo_to_access => ingress_fifo_to_access,
                                                ingress_fifo_address_from_read_ptr => ingress_fifo_address_from_read_ptr,
                                                ingress_fifo_event_type => ingress_fifo_event_type,

                                                ingress_sram_data_op => ingress_sram_data_op,
                                                ingress_sram_data_reg_hold => ingress_sram_data_reg_hold,
                                                ingress_sram_address_op => ingress_sram_address_op );

            io_ingress_fifos ingress_fifos( int_clock <- int_clock,
                                            int_reset <= int_reset,
                                            fifo_op <= ingress_fifo_op,
                                            fifo_op_to_status <= ingress_fifo_op_to_status,
                                            fifo_address_from_read_ptr <= ingress_fifo_address_from_read_ptr,
                                            fifo_address => ingress_fifo_address,
                                            fifo_event_type <= ingress_fifo_event_type,
                                            fifo_to_access <= ingress_fifo_to_access,

                                            status_fifo_empty => status_fifo_empty,
                                            status_fifo_full => status_fifo_full,
                                            status_fifo_overflowed => status_fifo_overflowed,
                                            status_fifo_underflowed => status_fifo_underflowed,

                                            rx_data_fifo_empty => rx_data_fifo_empty,
                                            rx_data_fifo_watermark => rx_data_fifo_watermark,
                                            rx_data_fifo_full => rx_data_fifo_full,
                                            rx_data_fifo_overflowed => rx_data_fifo_overflowed,
                                            rx_data_fifo_underflowed => rx_data_fifo_underflowed,

                                            event_from_status => ingress_event_from_status,
                                            event_fifo => ingress_event_fifo,
                                            event_empty => ingress_event_empty,
                                            event_watermark => ingress_event_watermark,

                                            cfg_base_address <= cfg_base_address,
                                            cfg_size_m_one <= cfg_size_m_one,
                                            cfg_watermark <= cfg_watermark,
                                            read_cfg_status => ingress_fifo_cfg_status );

        }

    /*b Ingress SRAM operation, data and address selectors
     */
    ingress_sram_controls "Ingress SRAM controls":
        {
            /*b Status timer
             */
            status_timer <= status_timer+1;

            if (!ingress_sram_data_reg_hold)
            {
                ingress_data_reg <= status_rx_data_fifo_data;
            }

            /*b Handle the data op
             */
            //   write timer value
            //   write ingress status data value
            //   write ingress rx data value
            //   ?write postbus data value
            //   read
            ingress_sram_write = 0;
            ingress_sram_read = 0;
            ingress_sram_write_data = ingress_data_reg;
            full_switch ( ingress_sram_data_op )
                {
                case io_sram_data_op_none:
                {
                    ingress_sram_write = 0;
                    ingress_sram_read = 0;
                    ingress_sram_write_data = ingress_data_reg;
                }
                case io_sram_data_op_write_time:
                {
                    ingress_sram_write = 1;
                    ingress_sram_write_data = status_timer;
                }
                case io_sram_data_op_write_data_reg:
                {
                    ingress_sram_write = 1;
                    ingress_sram_write_data = ingress_data_reg;
                }
                case io_sram_data_op_write_data:
                {
                    ingress_sram_write = 1;
                    ingress_sram_write_data = ingress_data_reg;
                }
                case io_sram_data_op_read:
                {
                    ingress_sram_read = 1;
                }
                case io_sram_data_op_read_fifo_status:
                {
                    ingress_sram_read = 0;
                }
                }


            /*b Handle the SRAM address
             */
            ingress_sram_address = ingress_fifo_address;
            full_switch ( ingress_sram_address_op )
                {
                case io_sram_address_op_egress_addressed:
                {
                    //ingress_sram_address = ingress_data_address;
                }
                case io_sram_address_op_postbus_addressed:
                {
                    //ingress_sram_address = ingress_postbus_address;
                }
                case io_sram_address_op_fifo_ptr:
                {
                    ingress_sram_address = ingress_fifo_address;
                }
                case io_sram_address_op_fifo_ptr_set_bit_0:
                {
                    ingress_sram_address = ingress_fifo_address;
                    ingress_sram_address[0] = 1;
                }
                }
        }

    /*b Ingress SRAM (RxData and status)
     */
    ingress_sram "Ingress sram":
        {
            memory_s_sp_2048_x_32 ingress_sram( sram_clock <- int_clock,
                                                sram_read <= ingress_sram_read,
                                                sram_write <= ingress_sram_write,
                                                sram_address <= ingress_sram_address,
                                                sram_write_data <= ingress_sram_write_data,
                                                sram_read_data => ingress_sram_read_data );
        }

    /*b IO cmd/tx data slot interface
     */
    io_cmd_tx_data_slot_interface "IO command and transmit data slot interface":
        {
            // note that the tx data interface runs at half speed, effectively, as a handled request will always be followed by an idle - this needs to be taken into account by the users
            io_slot_egr_data_ack = !tx_data_req; // if we do not have a request pending, then acknowledge anything if it arrives, coz we will make it pending
            if (tx_data_ack)
            {
                tx_data_req <= 0;
            }
            if (io_slot_egr_data_ack && io_slot_egr_data_req)
            {
                tx_data_req <= 1 ;
                tx_data_cmd <= io_slot_egr_data_cmd;
                tx_data_req_num <= io_slot_egr_data_slot;
            }
            last_io_slot_egr_cmd_ready <= io_slot_egr_cmd_ready;
            for (i; 4)
            {
                if ((!io_slot_egr_cmd_ready[i]) && (last_io_slot_egr_cmd_ready[i])) // on a cmd read the ready goes away - so our 'available' can clear to be filled again
                {
                    cmd_available_bus[i] <= 0;
                }
                if (cmd_valid && (i==cmd_valid_number)) // as soon as a read occurs though we need to set our indication, so that back-to-back commands to the same slot do not occur without a toggle from the I/O
                {
                    cmd_available_bus[i] <= 1;
                }
            }

            io_slot_egr_cmd_write <= 0;
            io_slot_egr_data_write <= 0;
            if (cmd_valid) 
            {
                io_slot_egr_slot <= cmd_valid_number;
                io_slot_egr_cmd_write <= 1;
                io_slot_egr_data <= egress_sram_read_data;
            }
            tx_data_read_being_presented <= tx_data_ack;
            tx_data_slot_being_presented <= tx_data_req_num;
            tx_data_reading              <= tx_data_read_being_presented;
            tx_data_slot_reading         <= tx_data_req_num;
            if (tx_data_reading)
            {
                io_slot_egr_slot <= tx_data_slot_reading;
                io_slot_egr_data_write <= 1;
                io_slot_egr_data <= egress_sram_read_data;
            }
        }

    /*b Command and TxData FIFO ptrs and their arbiter
     */
    comb bit[io_cmd_timestamp_length+2]io_timer;
    command_fifos_and_arbiter "Command, Tx data fifos, and arbiter":
        {
            io_timer = status_timer[io_cmd_timestamp_length+2;0];
            io_egress_control egress_control( int_clock <- int_clock,
                                              int_reset <= int_reset,

                                              io_timer <= io_timer,
                                              cmd_valid => cmd_valid,
                                              cmd_valid_number => cmd_valid_number,
                                              cmd_available <= cmd_available_bus,

                                              tx_data_req <= tx_data_req,
                                              tx_data_req_fifo <= tx_data_req_num,
                                              tx_data_ack => tx_data_ack,
                                              tx_data_cmd <= tx_data_cmd,

                                              postbus_req <= egress_postbus_req,
                                              postbus_ack => egress_postbus_ack,

                                              postbus_fifo_op <= egress_postbus_fifo_op,
                                              postbus_fifo_address_from_read_ptr <= egress_postbus_fifo_address_from_read_ptr,
                                              postbus_fifo_op_to_cmd <= egress_postbus_fifo_op_to_cmd_status,
                                              postbus_fifo_event_type <= egress_postbus_fifo_event_type,
                                              postbus_fifo_to_access <= egress_postbus_fifo_to_access,

                                              postbus_sram_data_op <= egress_postbus_sram_data_op,
                                              postbus_sram_address_op <= egress_postbus_sram_address_op,

                                              egress_fifo_op => egress_fifo_op,
                                              egress_fifo_op_to_cmd => egress_fifo_op_to_cmd,
                                              egress_fifo_to_access => egress_fifo_to_access,
                                              egress_fifo_address_from_read_ptr => egress_fifo_address_from_read_ptr,
                                              egress_fifo_event_type => egress_fifo_event_type,
                                              egress_cmd_fifo_empty <= cmd_fifo_empty,

                                              egress_sram_data_op => egress_sram_data_op,
                                              egress_sram_data_reg_op => egress_sram_data_reg_op,
                                              egress_sram_address_op => egress_sram_address_op,
                                              egress_sram_read_data <= egress_sram_read_data );

            io_egress_fifos egress_fifos( int_clock <- int_clock,
                                          int_reset <= int_reset,
                                          fifo_op <= egress_fifo_op,
                                          fifo_op_to_cmd <= egress_fifo_op_to_cmd,
                                          fifo_address_from_read_ptr <= egress_fifo_address_from_read_ptr,
                                          fifo_address => egress_fifo_address,
                                          fifo_event_type <= egress_fifo_event_type,
                                          fifo_to_access <= egress_fifo_to_access,

                                          cmd_fifo_empty => cmd_fifo_empty,
                                          cmd_fifo_full => cmd_fifo_full,
                                          cmd_fifo_overflowed => cmd_fifo_overflowed,
                                          cmd_fifo_underflowed => cmd_fifo_underflowed,

                                          tx_data_fifo_empty => tx_data_fifo_empty,
                                          tx_data_fifo_watermark => tx_data_fifo_watermark,
                                          tx_data_fifo_full => tx_data_fifo_full,
                                          tx_data_fifo_overflowed => tx_data_fifo_overflowed,
                                          tx_data_fifo_underflowed => tx_data_fifo_underflowed,

                                          event_from_cmd => egress_event_from_cmd,
                                          event_fifo => egress_event_fifo,
                                          event_empty => egress_event_empty,
                                          event_watermark => egress_event_watermark,

                                          cfg_base_address <= cfg_base_address,
                                          cfg_size_m_one <= cfg_size_m_one,
                                          cfg_watermark <= cfg_watermark,
                                          read_cfg_status => egress_fifo_cfg_status );

        }

    /*b Egress SRAM operation, data and address selectors
     */
    clocked bit[32] last_postbus_write_data=0;
    egress_sram_controls "Egress SRAM controls":
        {
            /*b Handle the data op
             */
            //   write from postbus
            //   ?read to postbus
            //   write from data reg
            //   read data
            //   read command time
            //   read command value
            egress_sram_write = 0;
            egress_sram_read = 0;
            egress_sram_write_data = egress_data_reg;
            last_postbus_write_data <= postbus_write_data;
            full_switch ( egress_sram_data_op )
                {
                case io_sram_data_op_none:
                {
                    egress_sram_write = 0;
                    egress_sram_read = 0;
                }
                case io_sram_data_op_read:
                {
                    egress_sram_read = 1;
                }
                case io_sram_data_op_write_time:
                case io_sram_data_op_write_data_reg:
                case io_sram_data_op_write_postbus:
                {
                    egress_sram_write = 1;
                    egress_sram_write_data = last_postbus_write_data;
                }
                case io_sram_data_op_read_fifo_status:
                {
                    egress_sram_read = 0;
                }
                }

            /*b Handle the data reg - DOES NOTHING! should select the appropriate interface, but we have just one at present
             */
            full_switch ( egress_sram_data_reg_op )
                {
                case io_sram_data_reg_op_hold:
                {
                    egress_data_reg <= egress_data_reg;
                }
                }

            /*b Handle the SRAM address
             */
            egress_sram_address = egress_fifo_address;
            full_switch ( egress_sram_address_op )
                {
                case io_sram_address_op_egress_addressed:
                {
                    //egress_sram_address = egress_data_address;
                }
                case io_sram_address_op_postbus_addressed:
                {
                    //egress_sram_address = egress_postbus_address;
                }
                case io_sram_address_op_fifo_ptr:
                {
                    egress_sram_address = egress_fifo_address;
                }
                case io_sram_address_op_fifo_ptr_set_bit_0:
                {
                    egress_sram_address = egress_fifo_address;
                    egress_sram_address[0] = 1;
                }
                }
        }

    /*b Egress SRAM (TxData and control)
     */
    egress_sram "Egress sram":
        {
            memory_s_sp_2048_x_32 egress_sram( sram_clock <- int_clock,
                                               sram_read <= egress_sram_read,
                                               sram_write <= egress_sram_write,
                                               sram_address <= egress_sram_address,
                                               sram_write_data <= egress_sram_write_data,
                                               sram_read_data => egress_sram_read_data );
        }

    /*b Baud rate generators
     */
    brg "Baud rate generators":
        {
            io_baud_rate_generator brg0 ( io_clock <- int_clock,
                                          io_reset <= int_reset,
                                          counter_enable <= brg0_counter_enable, // or allow for daisychaining or divide-by-input-enable
                                          counter_reset <= brg0_counter_reset, // or allow for synchronization
                                          baud_clock_enable => brg0_baud_enable,
                                          set_clock_config <= brg0_set_config,
                                          config_baud_addition_value <= cfg_baud_addition_value,
                                          config_baud_subtraction_value <= cfg_baud_subtraction_value
                );

            io_baud_rate_generator brg1 ( io_clock <- int_clock,
                                          io_reset <= int_reset,
                                          counter_enable <= brg1_counter_enable, // or allow for daisychaining or divide-by-input-enable
                                          counter_reset <= brg1_counter_reset, // or allow for synchronization
                                          baud_clock_enable => brg1_baud_enable,
                                          set_clock_config <= brg1_set_config,
                                          config_baud_addition_value <= cfg_baud_addition_value,
                                          config_baud_subtraction_value <= cfg_baud_subtraction_value
                );
        }

    /*b Postbus interface
     */
    postbus_interface "Postbus source and target":
        {
            io_postbus pst( int_clock <- int_clock,
                            int_reset <= int_reset,

                            postbus_src_type => postbus_src_type,
                            postbus_src_data => postbus_src_data,
                            postbus_src_ack <= postbus_src_ack,

                            postbus_tgt_type <= postbus_tgt_type,
                            postbus_tgt_data <= postbus_tgt_data,
                            postbus_tgt_ack => postbus_tgt_ack,

                            egress_req => egress_postbus_req,
                            egress_ack <= egress_postbus_ack,

                            egress_fifo_op => egress_postbus_fifo_op,
                            egress_fifo_op_to_cmd_status => egress_postbus_fifo_op_to_cmd_status,
                            egress_fifo_to_access => egress_postbus_fifo_to_access,
                            egress_fifo_event_type => egress_postbus_fifo_event_type,
                            egress_fifo_address_from_read_ptr => egress_postbus_fifo_address_from_read_ptr,

                            egress_sram_address_op => egress_postbus_sram_address_op,
                            egress_sram_data_op => egress_postbus_sram_data_op,

                            egress_event_from_cmd <= egress_event_from_cmd,
                            egress_event_fifo <= egress_event_fifo,
                            egress_event_empty <= egress_event_empty,
                            egress_event_watermark <= egress_event_watermark,

                            ingress_req => ingress_postbus_req,
                            ingress_ack <= ingress_postbus_ack,

                            ingress_fifo_op => ingress_postbus_fifo_op,
                            ingress_fifo_op_to_cmd_status => ingress_postbus_fifo_op_to_cmd_status,
                            ingress_fifo_to_access => ingress_postbus_fifo_to_access,
                            ingress_fifo_event_type => ingress_postbus_fifo_event_type,
                            ingress_fifo_address_from_read_ptr => ingress_postbus_fifo_address_from_read_ptr,

                            ingress_sram_address_op => ingress_postbus_sram_address_op,
                            ingress_sram_data_op => ingress_postbus_sram_data_op,

                            ingress_event_from_status <= ingress_event_from_status,
                            ingress_event_fifo <= ingress_event_fifo,
                            ingress_event_empty <= ingress_event_empty,
                            ingress_event_watermark <= ingress_event_watermark,

                            read_data <= postbus_src_read_data,

                            configuration_write => postbus_configuration_write,
                            write_address => postbus_write_address,
                            write_data => postbus_write_data );
            full_switch (postbus_src_read_data_source)
            {
            case postbus_src_read_data_source_ingress_fifo_status:
            case postbus_src_read_data_source_egress_fifo_status:
            {
                postbus_src_read_data = sram_read_data_fifo_status;
            }
            case postbus_src_read_data_source_ingress_sram:
            {
                postbus_src_read_data = ingress_sram_read_data; // if last but one ingress_req and was 
            }
            case postbus_src_read_data_source_egress_sram:
            {
                postbus_src_read_data = egress_sram_read_data;
            }
            }
            postbus_src_read_data_source <= next_postbus_src_read_data_source;
            next_postbus_src_read_data_source <= postbus_src_read_data_source_egress_sram;
            if (ingress_postbus_req)
            {
                next_postbus_src_read_data_source <= postbus_src_read_data_source_ingress_sram;
                if (ingress_postbus_sram_data_op==io_sram_data_op_read_fifo_status)
                {
                    next_postbus_src_read_data_source <= postbus_src_read_data_source_ingress_fifo_status;
                }
            }
            else
            {
                next_postbus_src_read_data_source <= postbus_src_read_data_source_egress_sram;
                if (egress_postbus_sram_data_op==io_sram_data_op_read_fifo_status)
                {
                    next_postbus_src_read_data_source <= postbus_src_read_data_source_egress_fifo_status;
                }
            }
            sram_read_data_fifo_status <= ingress_fifo_cfg_status;
            if (next_postbus_src_read_data_source==postbus_src_read_data_source_egress_fifo_status)
            {
                sram_read_data_fifo_status <= egress_fifo_cfg_status;
            }
        }

    /*b Configuration registers for postbus to handle later
     */
    config "Config data tie downs for now":
        {
            brg0_counter_enable = 1;
            brg0_counter_reset = 0;

            brg1_counter_enable = 1;
            brg1_counter_reset = 0;

            brg0_set_config = 0;
            brg1_set_config = 0;

            io_slot_cfg_write <= 0;
            if (postbus_configuration_write)
            {
                part_switch (postbus_write_address[3;0])
                {
                case 0:
                case 1:
                case 2:
                case 3:
                {
                    io_slot_cfg_write <= 1;
                    io_slot_cfg_slot <= postbus_write_address[2;0];
                    io_slot_cfg_data <= postbus_write_data[8;0];
                }
                case 4:
                {
                    brg0_set_config = 1;
                }
                case 5:
                {
                    brg1_set_config = 1;
                }
                }
            }

            cfg_baud_addition_value = postbus_write_data[io_baud_rate_divider_size;0];
            cfg_baud_subtraction_value = postbus_write_data[io_baud_rate_divider_size;16];

            cfg_size_m_one = 0;
            cfg_watermark  = 0;
            cfg_base_address                      = postbus_write_data[io_sram_log_size;0];
            cfg_size_m_one[io_sram_log_size-1;0]  = postbus_write_data[io_sram_log_size-1;io_sram_log_size];
            cfg_watermark[io_sram_log_size-1;0]   = postbus_write_data[io_sram_log_size-1;2*io_sram_log_size-1];
        }

    /*b -------------------- Done
     */
}
