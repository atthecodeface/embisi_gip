/*a Memory stage methods
 */
/*f c_gip_full::mem_comb
 */
void c_gip_full::mem_comb( t_gip_pipeline_results *results )
{
    /*b No need to do anything here as the actual combinatorials derive from the previous clock edge - see the clock funcion for that operation
     */
}

/*f c_gip_full::mem_preclock
 */
void c_gip_full::mem_preclock( void )
{

    /*b Copy current to next
     */
    memcpy( &pd->mem.next_state, &pd->mem.state, sizeof(pd->mem.state) );

    /*b Record input state
     */
    pd->mem.next_state.mem_rd = pd->alu.mem_rd;
    pd->mem.next_state.gip_mem_op = pd->alu.gip_mem_op;
    pd->mem.next_state.mem_data_in = pd->alu.mem_data_in;
    pd->mem.next_state.mem_address = pd->alu.mem_address;

}

/*f c_gip_full::mem_clock
 */
void c_gip_full::mem_clock( void )
{
    int offset_in_word;
    unsigned int data;
    unsigned int address;

    /*b Debug
     */
    if (pd->verbose)
    {
        printf( "\t**:MEM OP %d at %08x with %08x Rd %d/%02x\n",
                pd->mem.state.gip_mem_op,
                pd->mem.state.mem_address,
                pd->mem.state.mem_data_in,
                pd->mem.state.mem_rd.type,
                pd->mem.state.mem_rd.data.r );
    }

    /*b Perform a memory write if required
     */
    address = pd->mem.state.mem_address;
    switch (pd->mem.state.gip_mem_op)
    {
    case gip_mem_op_store_word:
        pd->memory->write_memory( address, pd->mem.state.mem_data_in, 0xf );
        break;
    case gip_mem_op_store_half:
        offset_in_word = address&0x2;
        address &= ~2;
        pd->memory->write_memory( address, pd->mem.state.mem_data_in<<(8*offset_in_word), 3<<offset_in_word );
        break;
    case gip_mem_op_store_byte:
        offset_in_word = address&0x3;
        address &= ~3;
        pd->memory->write_memory( address, pd->mem.state.mem_data_in<<(8*offset_in_word), 1<<offset_in_word );
        break;
    default:
        break;
    }

    /*b Copy next to current
     */
    memcpy( &pd->mem.state, &pd->mem.next_state, sizeof(pd->mem.state) );

    /*b Perform a memory read if required
     */
    address = pd->mem.state.mem_address;
    switch (pd->mem.state.gip_mem_op)
    {
    case gip_mem_op_load_word:
        pd->mem.mem_result = pd->memory->read_memory( address );
        break;
    case gip_mem_op_load_half:
        data = pd->memory->read_memory( address );
        offset_in_word = address&0x2;
        data >>= 8*offset_in_word;
        pd->mem.mem_result = data;
        break;
    case gip_mem_op_load_byte:
        data = pd->memory->read_memory( address );
        offset_in_word = address&0x3;
        data >>= 8*offset_in_word;
        pd->mem.mem_result = data;
        break;
    default:
        break;
    }
}

