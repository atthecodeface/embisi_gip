module barrel_shift_32
(
    select, in, out
);
input [4:0]select;
input [31:0]in;
output [31:0]out;

endmodule
